module cpu (clk, reset, DI, IRQ, NMI, RDY, AB, DO, WE);
input clk;
input reset;
input IRQ;
input NMI;
input RDY;
output WE;
input [7:0] DI;
output [15:0] AB;
output [7:0] DO;
wire vdd = 1'b1;
wire gnd = 1'b0;
BUFX4 BUFX4_1 ( .A(RDY), .Y(RDY_bF_buf8) );
BUFX4 BUFX4_2 ( .A(RDY), .Y(RDY_bF_buf7) );
BUFX4 BUFX4_3 ( .A(RDY), .Y(RDY_bF_buf6) );
BUFX4 BUFX4_4 ( .A(RDY), .Y(RDY_bF_buf5) );
BUFX4 BUFX4_5 ( .A(RDY), .Y(RDY_bF_buf4) );
BUFX4 BUFX4_6 ( .A(RDY), .Y(RDY_bF_buf3) );
BUFX4 BUFX4_7 ( .A(RDY), .Y(RDY_bF_buf2) );
BUFX4 BUFX4_8 ( .A(RDY), .Y(RDY_bF_buf1) );
BUFX4 BUFX4_9 ( .A(RDY), .Y(RDY_bF_buf0) );
BUFX4 BUFX4_10 ( .A(new_wire_28), .Y(_799__bF_buf4) );
BUFX4 BUFX4_11 ( .A(new_wire_28), .Y(_799__bF_buf3) );
BUFX4 BUFX4_12 ( .A(new_wire_28), .Y(_799__bF_buf2) );
BUFX4 BUFX4_13 ( .A(new_wire_28), .Y(_799__bF_buf1) );
BUFX4 BUFX4_14 ( .A(new_wire_29), .Y(_799__bF_buf0) );
BUFX4 BUFX4_15 ( .A(clk), .Y(clk_bF_buf11) );
BUFX4 BUFX4_16 ( .A(clk), .Y(clk_bF_buf10) );
BUFX4 BUFX4_17 ( .A(clk), .Y(clk_bF_buf9) );
BUFX4 BUFX4_18 ( .A(clk), .Y(clk_bF_buf8) );
BUFX4 BUFX4_19 ( .A(clk), .Y(clk_bF_buf7) );
BUFX4 BUFX4_20 ( .A(clk), .Y(clk_bF_buf6) );
BUFX4 BUFX4_21 ( .A(clk), .Y(clk_bF_buf5) );
BUFX4 BUFX4_22 ( .A(clk), .Y(clk_bF_buf4) );
BUFX4 BUFX4_23 ( .A(clk), .Y(clk_bF_buf3) );
BUFX4 BUFX4_24 ( .A(clk), .Y(clk_bF_buf2) );
BUFX4 BUFX4_25 ( .A(clk), .Y(clk_bF_buf1) );
BUFX4 BUFX4_26 ( .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_27 ( .A(_1101_), .Y(_1101__bF_buf3) );
BUFX4 BUFX4_28 ( .A(_1101_), .Y(_1101__bF_buf2) );
BUFX4 BUFX4_29 ( .A(_1101_), .Y(_1101__bF_buf1) );
BUFX4 BUFX4_30 ( .A(_1101_), .Y(_1101__bF_buf0) );
BUFX4 BUFX4_31 ( .A(new_wire_84), .Y(_849__bF_buf4) );
BUFX4 BUFX4_32 ( .A(new_wire_84), .Y(_849__bF_buf3) );
BUFX4 BUFX4_33 ( .A(new_wire_84), .Y(_849__bF_buf2) );
BUFX4 BUFX4_34 ( .A(new_wire_84), .Y(_849__bF_buf1) );
BUFX4 BUFX4_35 ( .A(new_wire_85), .Y(_849__bF_buf0) );
BUFX4 BUFX4_36 ( .A(new_wire_96), .Y(_825__bF_buf4) );
BUFX4 BUFX4_37 ( .A(new_wire_96), .Y(_825__bF_buf3) );
BUFX4 BUFX4_38 ( .A(new_wire_96), .Y(_825__bF_buf2) );
BUFX4 BUFX4_39 ( .A(new_wire_96), .Y(_825__bF_buf1) );
BUFX4 BUFX4_40 ( .A(new_wire_97), .Y(_825__bF_buf0) );
BUFX2 BUFX2_1 ( .A(_155_), .Y(_155__bF_buf3) );
BUFX2 BUFX2_2 ( .A(_155_), .Y(_155__bF_buf2) );
BUFX2 BUFX2_3 ( .A(_155_), .Y(_155__bF_buf1) );
BUFX2 BUFX2_4 ( .A(_155_), .Y(_155__bF_buf0) );
BUFX4 BUFX4_41 ( .A(new_wire_112), .Y(_822__bF_buf4) );
BUFX4 BUFX4_42 ( .A(new_wire_112), .Y(_822__bF_buf3) );
BUFX4 BUFX4_43 ( .A(new_wire_112), .Y(_822__bF_buf2) );
BUFX4 BUFX4_44 ( .A(new_wire_112), .Y(_822__bF_buf1) );
BUFX4 BUFX4_45 ( .A(new_wire_113), .Y(_822__bF_buf0) );
BUFX4 BUFX4_46 ( .A(_152_), .Y(_152__bF_buf3) );
BUFX4 BUFX4_47 ( .A(_152_), .Y(_152__bF_buf2) );
BUFX2 BUFX2_5 ( .A(_152_), .Y(_152__bF_buf1) );
BUFX2 BUFX2_6 ( .A(_152_), .Y(_152__bF_buf0) );
BUFX4 BUFX4_48 ( .A(new_wire_128), .Y(_795__bF_buf4) );
BUFX4 BUFX4_49 ( .A(new_wire_128), .Y(_795__bF_buf3) );
BUFX4 BUFX4_50 ( .A(new_wire_128), .Y(_795__bF_buf2) );
BUFX4 BUFX4_51 ( .A(new_wire_128), .Y(_795__bF_buf1) );
BUFX4 BUFX4_52 ( .A(new_wire_129), .Y(_795__bF_buf0) );
BUFX4 BUFX4_53 ( .A(new_wire_140), .Y(_651__bF_buf4) );
BUFX4 BUFX4_54 ( .A(new_wire_140), .Y(_651__bF_buf3) );
BUFX4 BUFX4_55 ( .A(new_wire_140), .Y(_651__bF_buf2) );
BUFX4 BUFX4_56 ( .A(new_wire_140), .Y(_651__bF_buf1) );
BUFX4 BUFX4_57 ( .A(new_wire_141), .Y(_651__bF_buf0) );
BUFX4 BUFX4_58 ( .A(new_wire_152), .Y(_1070__bF_buf4) );
BUFX4 BUFX4_59 ( .A(new_wire_152), .Y(_1070__bF_buf3) );
BUFX4 BUFX4_60 ( .A(new_wire_152), .Y(_1070__bF_buf2) );
BUFX4 BUFX4_61 ( .A(new_wire_152), .Y(_1070__bF_buf1) );
BUFX4 BUFX4_62 ( .A(new_wire_153), .Y(_1070__bF_buf0) );
BUFX2 BUFX2_7 ( .A(_830_), .Y(_830__bF_buf3) );
BUFX2 BUFX2_8 ( .A(_830_), .Y(_830__bF_buf2) );
BUFX2 BUFX2_9 ( .A(_830_), .Y(_830__bF_buf1) );
BUFX2 BUFX2_10 ( .A(_830_), .Y(_830__bF_buf0) );
BUFX4 BUFX4_63 ( .A(_1631_), .Y(_1631__bF_buf3) );
BUFX4 BUFX4_64 ( .A(_1631_), .Y(_1631__bF_buf2) );
BUFX4 BUFX4_65 ( .A(_1631_), .Y(_1631__bF_buf1) );
BUFX4 BUFX4_66 ( .A(_1631_), .Y(_1631__bF_buf0) );
BUFX4 BUFX4_67 ( .A(new_wire_174), .Y(_1017__bF_buf7) );
BUFX4 BUFX4_68 ( .A(new_wire_174), .Y(_1017__bF_buf6) );
BUFX4 BUFX4_69 ( .A(new_wire_174), .Y(_1017__bF_buf5) );
BUFX4 BUFX4_70 ( .A(new_wire_174), .Y(_1017__bF_buf4) );
BUFX4 BUFX4_71 ( .A(new_wire_175), .Y(_1017__bF_buf3) );
BUFX4 BUFX4_72 ( .A(new_wire_175), .Y(_1017__bF_buf2) );
BUFX4 BUFX4_73 ( .A(new_wire_175), .Y(_1017__bF_buf1) );
BUFX4 BUFX4_74 ( .A(new_wire_175), .Y(_1017__bF_buf0) );
BUFX4 BUFX4_75 ( .A(_859_), .Y(_859__bF_buf3) );
BUFX4 BUFX4_76 ( .A(_859_), .Y(_859__bF_buf2) );
BUFX2 BUFX2_11 ( .A(_859_), .Y(_859__bF_buf1) );
BUFX2 BUFX2_12 ( .A(_859_), .Y(_859__bF_buf0) );
BUFX4 BUFX4_77 ( .A(_148_), .Y(_148__bF_buf3) );
BUFX2 BUFX2_13 ( .A(_148_), .Y(_148__bF_buf2) );
BUFX2 BUFX2_14 ( .A(_148_), .Y(_148__bF_buf1) );
BUFX2 BUFX2_15 ( .A(_148_), .Y(_148__bF_buf0) );
BUFX4 BUFX4_78 ( .A(_815_), .Y(_815__bF_buf3) );
BUFX4 BUFX4_79 ( .A(_815_), .Y(_815__bF_buf2) );
BUFX4 BUFX4_80 ( .A(_815_), .Y(_815__bF_buf1) );
BUFX4 BUFX4_81 ( .A(_815_), .Y(_815__bF_buf0) );
BUFX4 BUFX4_82 ( .A(_812_), .Y(_812__bF_buf3) );
BUFX2 BUFX2_16 ( .A(_812_), .Y(_812__bF_buf2) );
BUFX4 BUFX4_83 ( .A(_812_), .Y(_812__bF_buf1) );
BUFX4 BUFX4_84 ( .A(_812_), .Y(_812__bF_buf0) );
BUFX4 BUFX4_85 ( .A(new_wire_219), .Y(_809__bF_buf4) );
BUFX4 BUFX4_86 ( .A(new_wire_219), .Y(_809__bF_buf3) );
BUFX4 BUFX4_87 ( .A(new_wire_219), .Y(_809__bF_buf2) );
BUFX4 BUFX4_88 ( .A(new_wire_219), .Y(_809__bF_buf1) );
BUFX4 BUFX4_89 ( .A(new_wire_220), .Y(_809__bF_buf0) );
INVX1 INVX1_1 ( .A(PC_13_), .Y(_787_) );
NAND2X1 NAND2X1_1 ( .A(new_wire_231), .B(new_wire_233), .Y(_788_) );
INVX2 INVX2_1 ( .A(_788_), .Y(_789_) );
INVX1 INVX1_2 ( .A(new_wire_237), .Y(_790_) );
NOR2X1 NOR2X1_1 ( .A(new_wire_239), .B(_790_), .Y(_791_) );
NAND2X1 NAND2X1_2 ( .A(new_wire_235), .B(_791_), .Y(_792_) );
INVX1 INVX1_3 ( .A(state_4_), .Y(_793_) );
NOR2X1 NOR2X1_2 ( .A(new_wire_243), .B(_793_), .Y(_794_) );
INVX8 INVX8_1 ( .A(new_wire_245), .Y(_795_) );
NOR2X1 NOR2X1_3 ( .A(new_wire_134), .B(new_wire_241), .Y(_796_) );
INVX1 INVX1_4 ( .A(new_wire_243), .Y(_797_) );
NOR2X1 NOR2X1_4 ( .A(state_4_), .B(_797_), .Y(_798_) );
INVX8 INVX8_2 ( .A(new_wire_251), .Y(_799_) );
INVX1 INVX1_5 ( .A(new_wire_231), .Y(_800_) );
NOR2X1 NOR2X1_5 ( .A(new_wire_233), .B(_800_), .Y(_801_) );
AND2X2 AND2X2_1 ( .A(new_wire_237), .B(new_wire_239), .Y(_802_) );
NAND2X1 NAND2X1_3 ( .A(new_wire_255), .B(_801_), .Y(_803_) );
INVX1 INVX1_6 ( .A(new_wire_239), .Y(_804_) );
NOR2X1 NOR2X1_6 ( .A(new_wire_237), .B(_804_), .Y(_805_) );
NAND2X1 NAND2X1_4 ( .A(_801_), .B(new_wire_257), .Y(_806_) );
AOI22X1 AOI22X1_1 ( .A(new_wire_134), .B(new_wire_36), .C(_803_), .D(_806_), .Y(_807_) );
NOR2X1 NOR2X1_7 ( .A(new_wire_249), .B(new_wire_259), .Y(_808_) );
OR2X2 OR2X2_1 ( .A(new_wire_243), .B(state_4_), .Y(_809_) );
NOR2X1 NOR2X1_8 ( .A(new_wire_231), .B(new_wire_233), .Y(_810_) );
NAND2X1 NAND2X1_5 ( .A(new_wire_265), .B(new_wire_255), .Y(_811_) );
NOR2X1 NOR2X1_9 ( .A(new_wire_243), .B(state_4_), .Y(_812_) );
INVX1 INVX1_7 ( .A(new_wire_233), .Y(_813_) );
NOR2X1 NOR2X1_10 ( .A(new_wire_231), .B(_813_), .Y(_814_) );
NAND3X1 NAND3X1_1 ( .A(new_wire_217), .B(_791_), .C(new_wire_267), .Y(_815_) );
OAI21X1 OAI21X1_1 ( .A(new_wire_223), .B(_811_), .C(new_wire_205), .Y(_816_) );
NAND3X1 NAND3X1_2 ( .A(new_wire_215), .B(new_wire_257), .C(new_wire_267), .Y(_817_) );
OAI21X1 OAI21X1_2 ( .A(new_wire_221), .B(new_wire_241), .C(new_wire_269), .Y(_818_) );
NOR2X1 NOR2X1_11 ( .A(_816_), .B(_818_), .Y(_819_) );
NAND2X1 NAND2X1_6 ( .A(new_wire_261), .B(new_wire_272), .Y(_820_) );
INVX1 INVX1_8 ( .A(new_wire_276), .Y(_821_) );
NAND3X1 NAND3X1_3 ( .A(new_wire_217), .B(new_wire_265), .C(new_wire_255), .Y(_822_) );
INVX1 INVX1_9 ( .A(IRQ), .Y(_823_) );
INVX8 INVX8_3 ( .A(NMI_edge), .Y(_824_) );
OAI21X1 OAI21X1_3 ( .A(I), .B(_823_), .C(new_wire_279), .Y(_825_) );
NOR2X1 NOR2X1_12 ( .A(new_wire_98), .B(new_wire_118), .Y(_826_) );
OAI21X1 OAI21X1_4 ( .A(_826_), .B(_821_), .C(PC_13_), .Y(_827_) );
INVX2 INVX2_2 ( .A(I), .Y(_828_) );
NAND2X1 NAND2X1_7 ( .A(_823_), .B(new_wire_279), .Y(_829_) );
OAI21X1 OAI21X1_5 ( .A(_828_), .B(NMI_edge), .C(_829_), .Y(_830_) );
NOR2X1 NOR2X1_13 ( .A(new_wire_118), .B(_830__bF_buf0), .Y(_831_) );
NAND2X1 NAND2X1_8 ( .A(ABH_5_), .B(_831_), .Y(_832_) );
NAND2X1 NAND2X1_9 ( .A(new_wire_237), .B(_804_), .Y(_833_) );
NOR2X1 NOR2X1_14 ( .A(_788_), .B(new_wire_283), .Y(_834_) );
NAND2X1 NAND2X1_10 ( .A(new_wire_245), .B(new_wire_285), .Y(_835_) );
NAND2X1 NAND2X1_11 ( .A(new_wire_232), .B(_813_), .Y(_836_) );
NAND2X1 NAND2X1_12 ( .A(new_wire_238), .B(new_wire_239), .Y(_837_) );
NOR2X1 NOR2X1_15 ( .A(_837_), .B(_836_), .Y(_838_) );
OAI21X1 OAI21X1_6 ( .A(new_wire_245), .B(new_wire_251), .C(new_wire_287), .Y(_839_) );
NAND2X1 NAND2X1_13 ( .A(new_wire_240), .B(_790_), .Y(_840_) );
NOR2X1 NOR2X1_16 ( .A(_836_), .B(_840_), .Y(_841_) );
OAI21X1 OAI21X1_7 ( .A(new_wire_245), .B(new_wire_251), .C(_841_), .Y(_842_) );
NAND3X1 NAND3X1_4 ( .A(_835_), .B(_839_), .C(_842_), .Y(_843_) );
INVX1 INVX1_10 ( .A(DIHOLD_5_), .Y(_844_) );
NAND2X1 NAND2X1_14 ( .A(new_wire_10), .B(DI[5]), .Y(_845_) );
OAI21X1 OAI21X1_8 ( .A(new_wire_10), .B(_844_), .C(_845_), .Y(DIMUX_5_) );
INVX2 INVX2_3 ( .A(new_wire_295), .Y(_846_) );
NAND3X1 NAND3X1_5 ( .A(new_wire_215), .B(new_wire_235), .C(_791_), .Y(_847_) );
NAND2X1 NAND2X1_15 ( .A(new_wire_234), .B(_800_), .Y(_848_) );
NOR3X1 NOR3X1_1 ( .A(new_wire_221), .B(new_wire_283), .C(_848_), .Y(_849_) );
NOR3X1 NOR3X1_2 ( .A(new_wire_221), .B(_840_), .C(_848_), .Y(_850_) );
AOI21X1 AOI21X1_1 ( .A(new_wire_90), .B(ABH_5_), .C(new_wire_302), .Y(_851_) );
OAI21X1 OAI21X1_9 ( .A(new_wire_298), .B(new_wire_300), .C(_851_), .Y(_852_) );
AOI21X1 AOI21X1_2 ( .A(new_wire_289), .B(new_wire_293), .C(_852_), .Y(_853_) );
NAND3X1 NAND3X1_6 ( .A(_832_), .B(_853_), .C(_827_), .Y(_854_) );
NAND3X1 NAND3X1_7 ( .A(PC_5_), .B(new_wire_261), .C(new_wire_272), .Y(_855_) );
NOR2X1 NOR2X1_17 ( .A(_840_), .B(_848_), .Y(_856_) );
AOI22X1 AOI22X1_2 ( .A(new_wire_211), .B(new_wire_305), .C(new_wire_295), .D(new_wire_86), .Y(_857_) );
NAND3X1 NAND3X1_8 ( .A(PC_5_), .B(new_wire_211), .C(new_wire_285), .Y(_858_) );
INVX8 INVX8_4 ( .A(new_wire_118), .Y(_859_) );
INVX2 INVX2_4 ( .A(PC_5_), .Y(_860_) );
NOR2X1 NOR2X1_18 ( .A(new_wire_307), .B(new_wire_102), .Y(_861_) );
INVX1 INVX1_11 ( .A(ABL_5_), .Y(_862_) );
NAND2X1 NAND2X1_16 ( .A(IRQ), .B(_828_), .Y(_863_) );
AOI21X1 AOI21X1_3 ( .A(new_wire_309), .B(new_wire_279), .C(_862_), .Y(_864_) );
OAI21X1 OAI21X1_10 ( .A(_864_), .B(_861_), .C(new_wire_195), .Y(_865_) );
NAND3X1 NAND3X1_9 ( .A(_858_), .B(_865_), .C(_857_), .Y(_866_) );
AOI21X1 AOI21X1_4 ( .A(new_wire_295), .B(new_wire_289), .C(_866_), .Y(_867_) );
NAND3X1 NAND3X1_10 ( .A(PC_4_), .B(new_wire_261), .C(new_wire_272), .Y(_868_) );
AOI21X1 AOI21X1_5 ( .A(new_wire_94), .B(new_wire_312), .C(new_wire_302), .Y(_869_) );
INVX4 INVX4_1 ( .A(new_wire_300), .Y(_870_) );
NAND2X1 NAND2X1_17 ( .A(PC_4_), .B(new_wire_315), .Y(_871_) );
INVX2 INVX2_5 ( .A(PC_4_), .Y(_872_) );
NOR2X1 NOR2X1_19 ( .A(new_wire_318), .B(new_wire_102), .Y(_873_) );
INVX1 INVX1_12 ( .A(ABL_4_), .Y(_874_) );
AOI21X1 AOI21X1_6 ( .A(new_wire_309), .B(new_wire_279), .C(_874_), .Y(_875_) );
OAI21X1 OAI21X1_11 ( .A(_875_), .B(_873_), .C(new_wire_195), .Y(_876_) );
NAND3X1 NAND3X1_11 ( .A(_876_), .B(_871_), .C(_869_), .Y(_877_) );
AOI21X1 AOI21X1_7 ( .A(new_wire_312), .B(new_wire_289), .C(_877_), .Y(_878_) );
AOI22X1 AOI22X1_3 ( .A(_867_), .B(_855_), .C(_868_), .D(_878_), .Y(_879_) );
NAND3X1 NAND3X1_12 ( .A(PC_7_), .B(new_wire_261), .C(new_wire_272), .Y(_880_) );
AOI22X1 AOI22X1_4 ( .A(new_wire_215), .B(new_wire_305), .C(new_wire_320), .D(new_wire_86), .Y(_881_) );
NAND3X1 NAND3X1_13 ( .A(PC_7_), .B(new_wire_211), .C(new_wire_285), .Y(_882_) );
INVX2 INVX2_6 ( .A(PC_7_), .Y(_883_) );
NOR2X1 NOR2X1_20 ( .A(new_wire_323), .B(new_wire_98), .Y(_884_) );
INVX1 INVX1_13 ( .A(ABL_7_), .Y(_885_) );
AOI21X1 AOI21X1_8 ( .A(new_wire_309), .B(new_wire_280), .C(_885_), .Y(_886_) );
OAI21X1 OAI21X1_12 ( .A(_886_), .B(_884_), .C(_859__bF_buf0), .Y(_887_) );
NAND3X1 NAND3X1_14 ( .A(_882_), .B(_887_), .C(_881_), .Y(_888_) );
AOI21X1 AOI21X1_9 ( .A(new_wire_320), .B(new_wire_289), .C(_888_), .Y(_889_) );
NAND3X1 NAND3X1_15 ( .A(PC_6_), .B(new_wire_262), .C(new_wire_273), .Y(_890_) );
AOI21X1 AOI21X1_10 ( .A(new_wire_86), .B(new_wire_325), .C(new_wire_302), .Y(_891_) );
NAND2X1 NAND2X1_18 ( .A(PC_6_), .B(new_wire_315), .Y(_892_) );
INVX2 INVX2_7 ( .A(PC_6_), .Y(_893_) );
NOR2X1 NOR2X1_21 ( .A(new_wire_328), .B(new_wire_98), .Y(_894_) );
INVX1 INVX1_14 ( .A(ABL_6_), .Y(_895_) );
AOI21X1 AOI21X1_11 ( .A(new_wire_309), .B(new_wire_280), .C(_895_), .Y(_896_) );
OAI21X1 OAI21X1_13 ( .A(_896_), .B(_894_), .C(_859__bF_buf0), .Y(_897_) );
NAND3X1 NAND3X1_16 ( .A(_897_), .B(_892_), .C(_891_), .Y(_898_) );
AOI21X1 AOI21X1_12 ( .A(new_wire_325), .B(new_wire_290), .C(_898_), .Y(_899_) );
AOI22X1 AOI22X1_5 ( .A(_889_), .B(_880_), .C(_890_), .D(_899_), .Y(_900_) );
NAND2X1 NAND2X1_19 ( .A(_879_), .B(_900_), .Y(_901_) );
NAND3X1 NAND3X1_17 ( .A(PC_0_), .B(new_wire_262), .C(new_wire_273), .Y(_902_) );
OAI21X1 OAI21X1_14 ( .A(new_wire_249), .B(new_wire_259), .C(new_wire_330), .Y(_903_) );
INVX2 INVX2_8 ( .A(new_wire_330), .Y(_904_) );
INVX2 INVX2_9 ( .A(PC_0_), .Y(_905_) );
OAI22X1 OAI22X1_1 ( .A(new_wire_333), .B(new_wire_300), .C(_904_), .D(new_wire_209), .Y(_906_) );
NAND2X1 NAND2X1_20 ( .A(ABL_0_), .B(new_wire_104), .Y(_907_) );
OAI21X1 OAI21X1_15 ( .A(new_wire_333), .B(new_wire_98), .C(_907_), .Y(_908_) );
AOI21X1 AOI21X1_13 ( .A(_859__bF_buf0), .B(_908_), .C(_906_), .Y(_909_) );
AND2X2 AND2X2_2 ( .A(_909_), .B(_903_), .Y(_910_) );
INVX1 INVX1_15 ( .A(_842_), .Y(_911_) );
XOR2X1 XOR2X1_1 ( .A(new_wire_335), .B(backwards), .Y(_912_) );
OAI22X1 OAI22X1_2 ( .A(new_wire_118), .B(new_wire_99), .C(_912_), .D(new_wire_207), .Y(_913_) );
NOR2X1 NOR2X1_22 ( .A(new_wire_238), .B(new_wire_240), .Y(_914_) );
NAND2X1 NAND2X1_21 ( .A(new_wire_337), .B(new_wire_267), .Y(_915_) );
NAND3X1 NAND3X1_18 ( .A(new_wire_235), .B(new_wire_215), .C(new_wire_257), .Y(_916_) );
OAI21X1 OAI21X1_16 ( .A(new_wire_221), .B(new_wire_339), .C(new_wire_341), .Y(_917_) );
NOR3X1 NOR3X1_3 ( .A(_917_), .B(_913_), .C(_911_), .Y(_918_) );
NAND2X1 NAND2X1_22 ( .A(new_wire_251), .B(new_wire_287), .Y(_919_) );
NOR2X1 NOR2X1_23 ( .A(new_wire_283), .B(_836_), .Y(_920_) );
INVX1 INVX1_16 ( .A(new_wire_343), .Y(_921_) );
OAI21X1 OAI21X1_17 ( .A(new_wire_222), .B(_921_), .C(_919_), .Y(_922_) );
NAND2X1 NAND2X1_23 ( .A(new_wire_265), .B(new_wire_337), .Y(_923_) );
INVX2 INVX2_10 ( .A(_923_), .Y(_924_) );
OAI21X1 OAI21X1_18 ( .A(new_wire_287), .B(_924_), .C(new_wire_213), .Y(_925_) );
OAI21X1 OAI21X1_19 ( .A(new_wire_244), .B(new_wire_241), .C(_925_), .Y(_926_) );
NOR2X1 NOR2X1_24 ( .A(_922_), .B(_926_), .Y(_927_) );
AOI22X1 AOI22X1_6 ( .A(_918_), .B(_927_), .C(_902_), .D(_910_), .Y(_928_) );
OAI21X1 OAI21X1_20 ( .A(new_wire_249), .B(new_wire_259), .C(new_wire_345), .Y(_929_) );
NAND3X1 NAND3X1_19 ( .A(PC_1_), .B(new_wire_262), .C(new_wire_273), .Y(_930_) );
INVX2 INVX2_11 ( .A(new_wire_345), .Y(_931_) );
OAI22X1 OAI22X1_3 ( .A(new_wire_347), .B(new_wire_209), .C(res), .D(new_wire_269), .Y(_932_) );
INVX2 INVX2_12 ( .A(PC_1_), .Y(_933_) );
NOR2X1 NOR2X1_25 ( .A(new_wire_349), .B(new_wire_300), .Y(_934_) );
NOR2X1 NOR2X1_26 ( .A(_934_), .B(_932_), .Y(_935_) );
NAND2X1 NAND2X1_24 ( .A(ABL_1_), .B(new_wire_104), .Y(_936_) );
OAI21X1 OAI21X1_21 ( .A(new_wire_349), .B(new_wire_104), .C(_936_), .Y(_937_) );
NAND2X1 NAND2X1_25 ( .A(new_wire_199), .B(_937_), .Y(_938_) );
AND2X2 AND2X2_3 ( .A(_935_), .B(_938_), .Y(_939_) );
NAND3X1 NAND3X1_20 ( .A(_929_), .B(_930_), .C(_939_), .Y(_940_) );
NAND3X1 NAND3X1_21 ( .A(PC_3_), .B(new_wire_262), .C(new_wire_273), .Y(_941_) );
AOI21X1 AOI21X1_14 ( .A(new_wire_94), .B(new_wire_351), .C(new_wire_302), .Y(_942_) );
NAND2X1 NAND2X1_26 ( .A(PC_3_), .B(new_wire_315), .Y(_943_) );
INVX2 INVX2_13 ( .A(PC_3_), .Y(_944_) );
NOR2X1 NOR2X1_27 ( .A(new_wire_354), .B(new_wire_102), .Y(_945_) );
INVX1 INVX1_17 ( .A(ABL_3_), .Y(_946_) );
AOI21X1 AOI21X1_15 ( .A(new_wire_310), .B(new_wire_280), .C(_946_), .Y(_947_) );
OAI21X1 OAI21X1_22 ( .A(_947_), .B(_945_), .C(new_wire_195), .Y(_948_) );
NAND3X1 NAND3X1_22 ( .A(_948_), .B(_943_), .C(_942_), .Y(_949_) );
AOI21X1 AOI21X1_16 ( .A(new_wire_351), .B(new_wire_290), .C(_949_), .Y(_950_) );
NAND3X1 NAND3X1_23 ( .A(PC_2_), .B(new_wire_263), .C(new_wire_274), .Y(_951_) );
NOR2X1 NOR2X1_28 ( .A(res), .B(new_wire_280), .Y(_952_) );
INVX1 INVX1_18 ( .A(_952_), .Y(_953_) );
AOI22X1 AOI22X1_7 ( .A(new_wire_94), .B(new_wire_356), .C(new_wire_303), .D(_953_), .Y(_954_) );
NAND2X1 NAND2X1_27 ( .A(PC_2_), .B(new_wire_315), .Y(_955_) );
INVX2 INVX2_14 ( .A(PC_2_), .Y(_956_) );
NOR2X1 NOR2X1_29 ( .A(new_wire_360), .B(new_wire_102), .Y(_957_) );
INVX1 INVX1_19 ( .A(ABL_2_), .Y(_958_) );
AOI21X1 AOI21X1_17 ( .A(new_wire_310), .B(new_wire_281), .C(_958_), .Y(_959_) );
OAI21X1 OAI21X1_23 ( .A(_959_), .B(_957_), .C(new_wire_195), .Y(_960_) );
NAND3X1 NAND3X1_24 ( .A(_955_), .B(_960_), .C(_954_), .Y(_961_) );
AOI21X1 AOI21X1_18 ( .A(new_wire_356), .B(new_wire_290), .C(_961_), .Y(_962_) );
AOI22X1 AOI22X1_8 ( .A(_950_), .B(_941_), .C(_951_), .D(_962_), .Y(_963_) );
NAND3X1 NAND3X1_25 ( .A(_940_), .B(_928_), .C(_963_), .Y(_964_) );
NAND3X1 NAND3X1_26 ( .A(PC_11_), .B(new_wire_263), .C(new_wire_274), .Y(_965_) );
INVX1 INVX1_20 ( .A(DIHOLD_3_), .Y(_966_) );
NAND2X1 NAND2X1_28 ( .A(new_wire_7), .B(DI[3]), .Y(_967_) );
OAI21X1 OAI21X1_24 ( .A(new_wire_7), .B(_966_), .C(_967_), .Y(DIMUX_3_) );
NAND3X1 NAND3X1_27 ( .A(new_wire_351), .B(new_wire_211), .C(new_wire_285), .Y(_968_) );
AOI21X1 AOI21X1_19 ( .A(new_wire_88), .B(ABH_3_), .C(new_wire_303), .Y(_969_) );
INVX1 INVX1_21 ( .A(ABH_3_), .Y(_970_) );
AOI21X1 AOI21X1_20 ( .A(new_wire_310), .B(new_wire_281), .C(_970_), .Y(_971_) );
INVX2 INVX2_15 ( .A(PC_11_), .Y(_972_) );
NOR2X1 NOR2X1_30 ( .A(new_wire_364), .B(new_wire_103), .Y(_973_) );
OAI21X1 OAI21X1_25 ( .A(_971_), .B(_973_), .C(new_wire_199), .Y(_974_) );
NAND3X1 NAND3X1_28 ( .A(_968_), .B(_974_), .C(_969_), .Y(_975_) );
AOI21X1 AOI21X1_21 ( .A(new_wire_290), .B(new_wire_362), .C(_975_), .Y(_976_) );
NAND3X1 NAND3X1_29 ( .A(PC_10_), .B(new_wire_263), .C(new_wire_274), .Y(_977_) );
MUX2X1 MUX2X1_1 ( .A(DI[2]), .B(DIHOLD_2_), .S(new_wire_10), .Y(_978_) );
INVX2 INVX2_16 ( .A(new_wire_366), .Y(DIMUX_2_) );
NAND2X1 NAND2X1_29 ( .A(new_wire_356), .B(new_wire_316), .Y(_979_) );
AOI21X1 AOI21X1_22 ( .A(new_wire_92), .B(ABH_2_), .C(new_wire_303), .Y(_980_) );
INVX1 INVX1_22 ( .A(ABH_2_), .Y(_981_) );
AOI21X1 AOI21X1_23 ( .A(new_wire_310), .B(new_wire_281), .C(_981_), .Y(_982_) );
INVX2 INVX2_17 ( .A(PC_10_), .Y(_983_) );
NOR2X1 NOR2X1_31 ( .A(new_wire_370), .B(new_wire_104), .Y(_984_) );
OAI21X1 OAI21X1_26 ( .A(_982_), .B(_984_), .C(new_wire_199), .Y(_985_) );
NAND3X1 NAND3X1_30 ( .A(_985_), .B(_979_), .C(_980_), .Y(_986_) );
AOI21X1 AOI21X1_24 ( .A(new_wire_291), .B(new_wire_368), .C(_986_), .Y(_987_) );
AOI22X1 AOI22X1_9 ( .A(_976_), .B(_965_), .C(_977_), .D(_987_), .Y(_988_) );
NAND3X1 NAND3X1_31 ( .A(PC_9_), .B(new_wire_263), .C(new_wire_274), .Y(_989_) );
INVX1 INVX1_23 ( .A(DIHOLD_1_), .Y(_990_) );
NAND2X1 NAND2X1_30 ( .A(new_wire_4), .B(DI[1]), .Y(_991_) );
OAI21X1 OAI21X1_27 ( .A(new_wire_4), .B(_990_), .C(_991_), .Y(DIMUX_1_) );
NAND3X1 NAND3X1_32 ( .A(new_wire_345), .B(new_wire_212), .C(new_wire_286), .Y(_992_) );
AOI21X1 AOI21X1_25 ( .A(new_wire_94), .B(ABH_1_), .C(new_wire_303), .Y(_993_) );
INVX1 INVX1_24 ( .A(ABH_1_), .Y(_994_) );
AOI21X1 AOI21X1_26 ( .A(new_wire_311), .B(new_wire_281), .C(_994_), .Y(_995_) );
INVX2 INVX2_18 ( .A(PC_9_), .Y(_996_) );
NOR2X1 NOR2X1_32 ( .A(_996_), .B(new_wire_103), .Y(_997_) );
OAI21X1 OAI21X1_28 ( .A(_995_), .B(_997_), .C(new_wire_196), .Y(_998_) );
NAND3X1 NAND3X1_33 ( .A(_992_), .B(_998_), .C(_993_), .Y(_999_) );
AOI21X1 AOI21X1_27 ( .A(new_wire_291), .B(new_wire_372), .C(_999_), .Y(_1000_) );
NAND3X1 NAND3X1_34 ( .A(PC_8_), .B(new_wire_264), .C(new_wire_275), .Y(_1001_) );
INVX1 INVX1_25 ( .A(DIHOLD_0_), .Y(_1002_) );
NAND2X1 NAND2X1_31 ( .A(new_wire_10), .B(DI[0]), .Y(_1003_) );
OAI21X1 OAI21X1_29 ( .A(new_wire_11), .B(_1002_), .C(_1003_), .Y(DIMUX_0_) );
NAND2X1 NAND2X1_32 ( .A(new_wire_330), .B(new_wire_316), .Y(_1004_) );
AOI21X1 AOI21X1_28 ( .A(new_wire_95), .B(ABH_0_), .C(new_wire_304), .Y(_1005_) );
INVX1 INVX1_26 ( .A(ABH_0_), .Y(_1006_) );
AOI21X1 AOI21X1_29 ( .A(new_wire_311), .B(new_wire_282), .C(_1006_), .Y(_1007_) );
INVX2 INVX2_19 ( .A(PC_8_), .Y(_1008_) );
NOR2X1 NOR2X1_33 ( .A(_1008_), .B(new_wire_105), .Y(_1009_) );
OAI21X1 OAI21X1_30 ( .A(_1007_), .B(_1009_), .C(new_wire_199), .Y(_1010_) );
NAND3X1 NAND3X1_35 ( .A(_1010_), .B(_1004_), .C(_1005_), .Y(_1011_) );
AOI21X1 AOI21X1_30 ( .A(new_wire_291), .B(new_wire_374), .C(_1011_), .Y(_1012_) );
AOI22X1 AOI22X1_10 ( .A(_1000_), .B(_989_), .C(_1001_), .D(_1012_), .Y(_1013_) );
NAND2X1 NAND2X1_33 ( .A(_988_), .B(_1013_), .Y(_1014_) );
NOR3X1 NOR3X1_4 ( .A(_901_), .B(_1014_), .C(_964_), .Y(_1015_) );
INVX2 INVX2_20 ( .A(PC_12_), .Y(_1016_) );
INVX8 INVX8_5 ( .A(new_wire_19), .Y(_1017_) );
OR2X2 OR2X2_2 ( .A(new_wire_11), .B(DIHOLD_4_), .Y(_1018_) );
OAI21X1 OAI21X1_31 ( .A(new_wire_185), .B(DI[4]), .C(_1018_), .Y(_1019_) );
INVX2 INVX2_21 ( .A(new_wire_378), .Y(DIMUX_4_) );
INVX2 INVX2_22 ( .A(ABH_4_), .Y(_1020_) );
OAI21X1 OAI21X1_32 ( .A(_1020_), .B(new_wire_209), .C(new_wire_269), .Y(_1021_) );
AOI21X1 AOI21X1_31 ( .A(new_wire_312), .B(new_wire_316), .C(_1021_), .Y(_1022_) );
NOR2X1 NOR2X1_34 ( .A(new_wire_376), .B(new_wire_105), .Y(_1023_) );
NOR2X1 NOR2X1_35 ( .A(_1020_), .B(_830__bF_buf0), .Y(_1024_) );
OAI21X1 OAI21X1_33 ( .A(_1023_), .B(_1024_), .C(new_wire_200), .Y(_1025_) );
NAND2X1 NAND2X1_34 ( .A(_1025_), .B(_1022_), .Y(_1026_) );
AOI21X1 AOI21X1_32 ( .A(new_wire_291), .B(DIMUX_4_), .C(_1026_), .Y(_1027_) );
OAI21X1 OAI21X1_34 ( .A(new_wire_376), .B(new_wire_276), .C(_1027_), .Y(_1028_) );
AOI21X1 AOI21X1_33 ( .A(_1015_), .B(new_wire_380), .C(_854_), .Y(_1029_) );
AND2X2 AND2X2_4 ( .A(_879_), .B(_900_), .Y(_1030_) );
NAND2X1 NAND2X1_35 ( .A(_940_), .B(_928_), .Y(_1031_) );
INVX1 INVX1_27 ( .A(_941_), .Y(_1032_) );
OAI21X1 OAI21X1_35 ( .A(new_wire_249), .B(new_wire_259), .C(new_wire_351), .Y(_1033_) );
AND2X2 AND2X2_5 ( .A(_942_), .B(_943_), .Y(_1034_) );
NAND3X1 NAND3X1_36 ( .A(_1033_), .B(_948_), .C(_1034_), .Y(_1035_) );
INVX1 INVX1_28 ( .A(_951_), .Y(_1036_) );
OAI21X1 OAI21X1_36 ( .A(new_wire_250), .B(new_wire_260), .C(new_wire_356), .Y(_1037_) );
AND2X2 AND2X2_6 ( .A(_954_), .B(_955_), .Y(_1038_) );
NAND3X1 NAND3X1_37 ( .A(_1037_), .B(_960_), .C(_1038_), .Y(_1039_) );
OAI22X1 OAI22X1_4 ( .A(_1035_), .B(_1032_), .C(_1036_), .D(_1039_), .Y(_1040_) );
NOR2X1 NOR2X1_36 ( .A(_1040_), .B(_1031_), .Y(_1041_) );
AND2X2 AND2X2_7 ( .A(_988_), .B(_1013_), .Y(_1042_) );
NAND3X1 NAND3X1_38 ( .A(_1030_), .B(_1042_), .C(_1041_), .Y(_1043_) );
NAND2X1 NAND2X1_36 ( .A(new_wire_380), .B(_854_), .Y(_1044_) );
OAI21X1 OAI21X1_37 ( .A(_1044_), .B(_1043_), .C(new_wire_16), .Y(_1045_) );
OAI22X1 OAI22X1_5 ( .A(_787_), .B(new_wire_11), .C(_1029_), .D(_1045_), .Y(_9__13_) );
NAND2X1 NAND2X1_37 ( .A(PC_14_), .B(new_wire_185), .Y(_1046_) );
NOR2X1 NOR2X1_37 ( .A(_1044_), .B(_1043_), .Y(_1047_) );
OAI21X1 OAI21X1_38 ( .A(_826_), .B(_821_), .C(PC_14_), .Y(_1048_) );
INVX1 INVX1_29 ( .A(ABH_6_), .Y(_1049_) );
OAI21X1 OAI21X1_39 ( .A(_1049_), .B(new_wire_209), .C(new_wire_269), .Y(_1050_) );
AOI21X1 AOI21X1_34 ( .A(new_wire_325), .B(new_wire_316), .C(_1050_), .Y(_1051_) );
MUX2X1 MUX2X1_2 ( .A(DI[6]), .B(DIHOLD_6_), .S(new_wire_25), .Y(_1052_) );
INVX2 INVX2_23 ( .A(new_wire_382), .Y(DIMUX_6_) );
AOI22X1 AOI22X1_11 ( .A(ABH_6_), .B(_831_), .C(new_wire_384), .D(new_wire_292), .Y(_1053_) );
NAND3X1 NAND3X1_39 ( .A(_1051_), .B(_1053_), .C(_1048_), .Y(_1054_) );
NOR2X1 NOR2X1_38 ( .A(_1054_), .B(_1047_), .Y(_1055_) );
AND2X2 AND2X2_8 ( .A(_854_), .B(new_wire_380), .Y(_1056_) );
NAND3X1 NAND3X1_40 ( .A(_1056_), .B(_1054_), .C(_1015_), .Y(_1057_) );
NAND2X1 NAND2X1_38 ( .A(new_wire_16), .B(_1057_), .Y(_1058_) );
OAI21X1 OAI21X1_40 ( .A(_1058_), .B(_1055_), .C(_1046_), .Y(_9__14_) );
INVX1 INVX1_30 ( .A(PC_15_), .Y(_1059_) );
OAI21X1 OAI21X1_41 ( .A(_826_), .B(_821_), .C(PC_15_), .Y(_1060_) );
INVX1 INVX1_31 ( .A(ABH_7_), .Y(_1061_) );
OAI21X1 OAI21X1_42 ( .A(_1061_), .B(new_wire_210), .C(new_wire_270), .Y(_1062_) );
AOI21X1 AOI21X1_35 ( .A(ABH_7_), .B(_831_), .C(_1062_), .Y(_1063_) );
MUX2X1 MUX2X1_3 ( .A(DI[7]), .B(DIHOLD_7_), .S(new_wire_11), .Y(_1064_) );
INVX2 INVX2_24 ( .A(new_wire_386), .Y(DIMUX_7_) );
AOI22X1 AOI22X1_12 ( .A(new_wire_320), .B(new_wire_317), .C(new_wire_388), .D(new_wire_292), .Y(_1065_) );
NAND3X1 NAND3X1_41 ( .A(_1063_), .B(_1065_), .C(_1060_), .Y(_1066_) );
INVX1 INVX1_32 ( .A(_1066_), .Y(_1067_) );
NAND3X1 NAND3X1_42 ( .A(_1054_), .B(_1067_), .C(_1047_), .Y(_1068_) );
AOI21X1 AOI21X1_36 ( .A(_1057_), .B(_1066_), .C(new_wire_185), .Y(_1069_) );
AOI22X1 AOI22X1_13 ( .A(new_wire_185), .B(_1059_), .C(_1068_), .D(_1069_), .Y(_9__15_) );
NOR2X1 NOR2X1_39 ( .A(new_wire_187), .B(new_wire_122), .Y(_1070_) );
NAND2X1 NAND2X1_39 ( .A(new_wire_337), .B(_801_), .Y(_1071_) );
NOR2X1 NOR2X1_40 ( .A(new_wire_38), .B(new_wire_390), .Y(_1072_) );
INVX4 INVX4_2 ( .A(new_wire_394), .Y(_1073_) );
INVX1 INVX1_33 ( .A(IRHOLD_3_), .Y(_1074_) );
NAND2X1 NAND2X1_40 ( .A(new_wire_397), .B(new_wire_362), .Y(_1075_) );
OAI21X1 OAI21X1_43 ( .A(new_wire_397), .B(_1074_), .C(_1075_), .Y(_1076_) );
NAND2X1 NAND2X1_41 ( .A(new_wire_164), .B(_1076_), .Y(_1077_) );
NAND2X1 NAND2X1_42 ( .A(new_wire_394), .B(IRHOLD_2_), .Y(_1078_) );
OAI21X1 OAI21X1_44 ( .A(new_wire_394), .B(new_wire_366), .C(_1078_), .Y(_1079_) );
AND2X2 AND2X2_9 ( .A(_1079_), .B(new_wire_164), .Y(_1080_) );
NOR2X1 NOR2X1_41 ( .A(new_wire_399), .B(_1077_), .Y(_1081_) );
MUX2X1 MUX2X1_4 ( .A(new_wire_372), .B(IRHOLD_1_), .S(new_wire_397), .Y(_1082_) );
NOR2X1 NOR2X1_42 ( .A(new_wire_100), .B(_1082_), .Y(_1083_) );
MUX2X1 MUX2X1_5 ( .A(new_wire_374), .B(IRHOLD_0_), .S(new_wire_397), .Y(_1084_) );
NOR2X1 NOR2X1_43 ( .A(new_wire_100), .B(new_wire_401), .Y(_1085_) );
NOR2X1 NOR2X1_44 ( .A(_1083_), .B(_1085_), .Y(_1086_) );
NAND2X1 NAND2X1_43 ( .A(new_wire_403), .B(_1081_), .Y(_1087_) );
NAND2X1 NAND2X1_44 ( .A(new_wire_394), .B(IRHOLD_7_), .Y(_1088_) );
OAI21X1 OAI21X1_45 ( .A(new_wire_395), .B(new_wire_386), .C(_1088_), .Y(_1089_) );
NAND2X1 NAND2X1_45 ( .A(_830__bF_buf0), .B(_1089_), .Y(_1090_) );
NAND2X1 NAND2X1_46 ( .A(new_wire_395), .B(IRHOLD_4_), .Y(_1091_) );
OAI21X1 OAI21X1_46 ( .A(new_wire_395), .B(new_wire_378), .C(_1091_), .Y(_1092_) );
MUX2X1 MUX2X1_6 ( .A(new_wire_293), .B(IRHOLD_5_), .S(new_wire_398), .Y(_1093_) );
NOR2X1 NOR2X1_45 ( .A(new_wire_106), .B(new_wire_413), .Y(_1094_) );
AOI21X1 AOI21X1_37 ( .A(_830__bF_buf2), .B(new_wire_411), .C(new_wire_415), .Y(_1095_) );
NAND2X1 NAND2X1_47 ( .A(new_wire_407), .B(_1095_), .Y(_1096_) );
NOR2X1 NOR2X1_46 ( .A(_1096_), .B(new_wire_405), .Y(_1097_) );
AOI22X1 AOI22X1_14 ( .A(new_wire_176), .B(new_wire_392), .C(new_wire_156), .D(_1097_), .Y(_1098_) );
NOR2X1 NOR2X1_47 ( .A(new_wire_229), .B(_921_), .Y(_1099_) );
INVX4 INVX4_3 ( .A(_1099_), .Y(_1100_) );
INVX8 INVX8_6 ( .A(new_wire_160), .Y(_1101_) );
AND2X2 AND2X2_10 ( .A(new_wire_411), .B(_830__bF_buf2), .Y(_1102_) );
OAI21X1 OAI21X1_47 ( .A(_1079_), .B(_1076_), .C(new_wire_164), .Y(_1103_) );
NAND3X1 NAND3X1_43 ( .A(new_wire_421), .B(_1103_), .C(new_wire_403), .Y(_1104_) );
OAI22X1 OAI22X1_6 ( .A(new_wire_22), .B(new_wire_418), .C(new_wire_76), .D(_1104_), .Y(_1105_) );
INVX1 INVX1_34 ( .A(new_wire_337), .Y(_1106_) );
NOR2X1 NOR2X1_48 ( .A(_836_), .B(_1106_), .Y(_1107_) );
NOR2X1 NOR2X1_49 ( .A(_797_), .B(_793_), .Y(_1108_) );
NAND2X1 NAND2X1_48 ( .A(_1108_), .B(_1107_), .Y(_1109_) );
NAND3X1 NAND3X1_44 ( .A(new_wire_265), .B(new_wire_338), .C(_1108_), .Y(_1110_) );
INVX1 INVX1_35 ( .A(_1110_), .Y(_1111_) );
NAND2X1 NAND2X1_49 ( .A(new_wire_13), .B(_1111_), .Y(_1112_) );
OAI21X1 OAI21X1_48 ( .A(new_wire_13), .B(_1109_), .C(_1112_), .Y(_1113_) );
NAND2X1 NAND2X1_50 ( .A(new_wire_246), .B(_1107_), .Y(_1114_) );
NAND2X1 NAND2X1_51 ( .A(new_wire_246), .B(_924_), .Y(_1115_) );
MUX2X1 MUX2X1_7 ( .A(_1114_), .B(_1115_), .S(new_wire_193), .Y(_1116_) );
NOR2X1 NOR2X1_50 ( .A(_1116_), .B(_1113_), .Y(_1117_) );
OAI21X1 OAI21X1_49 ( .A(new_wire_36), .B(_806_), .C(new_wire_193), .Y(_1118_) );
NAND2X1 NAND2X1_52 ( .A(new_wire_266), .B(new_wire_257), .Y(_1119_) );
OAI21X1 OAI21X1_50 ( .A(new_wire_36), .B(new_wire_425), .C(new_wire_19), .Y(_1120_) );
AND2X2 AND2X2_11 ( .A(_1118_), .B(_1120_), .Y(_1121_) );
NAND2X1 NAND2X1_53 ( .A(new_wire_213), .B(_841_), .Y(_1122_) );
NOR2X1 NOR2X1_51 ( .A(new_wire_223), .B(new_wire_425), .Y(_1123_) );
NAND2X1 NAND2X1_54 ( .A(new_wire_1), .B(_1123_), .Y(_1124_) );
OAI21X1 OAI21X1_51 ( .A(new_wire_13), .B(_1122_), .C(_1124_), .Y(_1125_) );
NOR2X1 NOR2X1_52 ( .A(_1121_), .B(_1125_), .Y(_1126_) );
NOR2X1 NOR2X1_53 ( .A(new_wire_134), .B(new_wire_425), .Y(_1127_) );
OAI21X1 OAI21X1_52 ( .A(new_wire_134), .B(_806_), .C(new_wire_193), .Y(_1128_) );
OAI21X1 OAI21X1_53 ( .A(new_wire_193), .B(_1127_), .C(_1128_), .Y(_1129_) );
NOR2X1 NOR2X1_54 ( .A(new_wire_229), .B(new_wire_390), .Y(_1130_) );
OAI21X1 OAI21X1_54 ( .A(new_wire_229), .B(_923_), .C(new_wire_13), .Y(_1131_) );
OAI21X1 OAI21X1_55 ( .A(new_wire_14), .B(_1130_), .C(_1131_), .Y(_1132_) );
AND2X2 AND2X2_12 ( .A(_1129_), .B(_1132_), .Y(_1133_) );
NAND3X1 NAND3X1_45 ( .A(_1133_), .B(_1117_), .C(_1126_), .Y(_1134_) );
NOR2X1 NOR2X1_55 ( .A(_1134_), .B(_1105_), .Y(_1135_) );
OAI21X1 OAI21X1_56 ( .A(new_wire_411), .B(_1076_), .C(_830__bF_buf2), .Y(_1136_) );
NOR2X1 NOR2X1_56 ( .A(_788_), .B(_837_), .Y(_1137_) );
INVX2 INVX2_25 ( .A(_1137_), .Y(_1138_) );
NOR2X1 NOR2X1_57 ( .A(new_wire_34), .B(new_wire_427), .Y(_1139_) );
NAND2X1 NAND2X1_55 ( .A(new_wire_164), .B(_1079_), .Y(_1140_) );
NOR2X1 NOR2X1_58 ( .A(new_wire_429), .B(new_wire_80), .Y(_1141_) );
AOI22X1 AOI22X1_15 ( .A(new_wire_176), .B(_1139_), .C(_1136_), .D(_1141_), .Y(_1142_) );
NAND2X1 NAND2X1_56 ( .A(new_wire_213), .B(_1137_), .Y(_1143_) );
INVX1 INVX1_36 ( .A(_1143_), .Y(_1144_) );
NAND2X1 NAND2X1_57 ( .A(new_wire_255), .B(new_wire_267), .Y(_1145_) );
OAI21X1 OAI21X1_57 ( .A(new_wire_227), .B(new_wire_431), .C(new_wire_1), .Y(_1146_) );
OAI21X1 OAI21X1_58 ( .A(new_wire_1), .B(_1144_), .C(_1146_), .Y(_1147_) );
NAND2X1 NAND2X1_58 ( .A(_1147_), .B(_1142_), .Y(_1148_) );
NOR2X1 NOR2X1_59 ( .A(new_wire_283), .B(_848_), .Y(_1149_) );
NAND2X1 NAND2X1_59 ( .A(new_wire_246), .B(_1149_), .Y(_1150_) );
NAND2X1 NAND2X1_60 ( .A(new_wire_19), .B(_1150_), .Y(_1151_) );
OAI21X1 OAI21X1_59 ( .A(new_wire_19), .B(new_wire_250), .C(_1151_), .Y(_1152_) );
INVX1 INVX1_37 ( .A(_1152_), .Y(_1153_) );
NAND2X1 NAND2X1_61 ( .A(new_wire_252), .B(_1149_), .Y(_1154_) );
NOR2X1 NOR2X1_60 ( .A(new_wire_38), .B(new_wire_241), .Y(_1155_) );
NAND2X1 NAND2X1_62 ( .A(new_wire_189), .B(new_wire_434), .Y(_1156_) );
OAI21X1 OAI21X1_60 ( .A(new_wire_189), .B(_1154_), .C(_1156_), .Y(_1157_) );
OR2X2 OR2X2_3 ( .A(_1153_), .B(_1157_), .Y(_1158_) );
NOR2X1 NOR2X1_61 ( .A(_1148_), .B(_1158_), .Y(_1159_) );
NAND2X1 NAND2X1_63 ( .A(new_wire_252), .B(new_wire_305), .Y(_1160_) );
NAND2X1 NAND2X1_64 ( .A(new_wire_235), .B(new_wire_258), .Y(_1161_) );
NOR2X1 NOR2X1_62 ( .A(new_wire_36), .B(new_wire_436), .Y(_1162_) );
NAND2X1 NAND2X1_65 ( .A(new_wire_194), .B(_1162_), .Y(_1163_) );
OAI21X1 OAI21X1_61 ( .A(new_wire_194), .B(_1160_), .C(_1163_), .Y(_1164_) );
MUX2X1 MUX2X1_8 ( .A(new_wire_270), .B(new_wire_341), .S(new_wire_14), .Y(_1165_) );
OR2X2 OR2X2_4 ( .A(_1164_), .B(_1165_), .Y(_1166_) );
NAND2X1 NAND2X1_66 ( .A(new_wire_4), .B(_912_), .Y(_1167_) );
OAI22X1 OAI22X1_7 ( .A(new_wire_4), .B(new_wire_301), .C(new_wire_207), .D(_1167_), .Y(_1168_) );
INVX1 INVX1_38 ( .A(_1168_), .Y(_1169_) );
NOR2X1 NOR2X1_63 ( .A(new_wire_138), .B(new_wire_436), .Y(_1170_) );
NAND2X1 NAND2X1_67 ( .A(new_wire_258), .B(new_wire_268), .Y(_1171_) );
OAI21X1 OAI21X1_62 ( .A(new_wire_138), .B(new_wire_438), .C(new_wire_20), .Y(_1172_) );
OAI21X1 OAI21X1_63 ( .A(new_wire_20), .B(_1170_), .C(_1172_), .Y(_1173_) );
NAND2X1 NAND2X1_68 ( .A(_1173_), .B(_1169_), .Y(_1174_) );
NOR2X1 NOR2X1_64 ( .A(_1174_), .B(_1166_), .Y(_1176_) );
NAND2X1 NAND2X1_69 ( .A(_1176_), .B(_1159_), .Y(_1177_) );
NAND2X1 NAND2X1_70 ( .A(_830__bF_buf1), .B(new_wire_411), .Y(_1178_) );
INVX2 INVX2_26 ( .A(new_wire_362), .Y(_1179_) );
OAI21X1 OAI21X1_64 ( .A(new_wire_398), .B(IRHOLD_3_), .C(_830__bF_buf0), .Y(_1180_) );
AOI21X1 AOI21X1_38 ( .A(new_wire_398), .B(_1179_), .C(_1180_), .Y(_1181_) );
NAND2X1 NAND2X1_71 ( .A(new_wire_429), .B(_1181_), .Y(_1182_) );
OAI21X1 OAI21X1_65 ( .A(new_wire_100), .B(_1082_), .C(_1085_), .Y(_1183_) );
NOR2X1 NOR2X1_65 ( .A(new_wire_445), .B(new_wire_443), .Y(_1184_) );
NAND2X1 NAND2X1_72 ( .A(new_wire_440), .B(_1184_), .Y(_1185_) );
NAND2X1 NAND2X1_73 ( .A(new_wire_429), .B(_1077_), .Y(_1186_) );
NOR2X1 NOR2X1_66 ( .A(new_wire_407), .B(new_wire_421), .Y(_1187_) );
OAI21X1 OAI21X1_66 ( .A(new_wire_100), .B(new_wire_401), .C(_1187_), .Y(_1188_) );
OAI21X1 OAI21X1_67 ( .A(_1186_), .B(_1188_), .C(_1185_), .Y(_1189_) );
OAI21X1 OAI21X1_68 ( .A(new_wire_343), .B(_1107_), .C(new_wire_246), .Y(_1190_) );
INVX1 INVX1_39 ( .A(new_wire_431), .Y(_1191_) );
NAND2X1 NAND2X1_74 ( .A(new_wire_252), .B(_1191_), .Y(_1192_) );
NAND3X1 NAND3X1_46 ( .A(_839_), .B(_1190_), .C(new_wire_447), .Y(_1193_) );
OAI21X1 OAI21X1_69 ( .A(new_wire_229), .B(new_wire_390), .C(_1109_), .Y(_1194_) );
NAND2X1 NAND2X1_75 ( .A(_800_), .B(_813_), .Y(_1195_) );
NOR2X1 NOR2X1_67 ( .A(new_wire_284), .B(_1195_), .Y(_1196_) );
NAND2X1 NAND2X1_76 ( .A(new_wire_217), .B(new_wire_449), .Y(_1197_) );
OAI21X1 OAI21X1_70 ( .A(new_wire_38), .B(new_wire_427), .C(_1197_), .Y(_1198_) );
NOR2X1 NOR2X1_68 ( .A(_1198_), .B(_1194_), .Y(_1199_) );
NAND3X1 NAND3X1_47 ( .A(new_wire_1), .B(_1193_), .C(_1199_), .Y(_1200_) );
NAND3X1 NAND3X1_48 ( .A(new_wire_256), .B(new_wire_266), .C(new_wire_252), .Y(_1201_) );
INVX1 INVX1_40 ( .A(_1201_), .Y(_1202_) );
NAND2X1 NAND2X1_77 ( .A(new_wire_5), .B(_1202_), .Y(_1203_) );
OAI21X1 OAI21X1_71 ( .A(new_wire_5), .B(_919_), .C(_1203_), .Y(_1204_) );
NAND2X1 NAND2X1_78 ( .A(new_wire_217), .B(new_wire_287), .Y(_1205_) );
NAND2X1 NAND2X1_79 ( .A(new_wire_247), .B(new_wire_449), .Y(_1206_) );
NOR2X1 NOR2X1_69 ( .A(store), .B(new_wire_335), .Y(_1207_) );
NAND2X1 NAND2X1_80 ( .A(new_wire_25), .B(_1207_), .Y(_1208_) );
OAI22X1 OAI22X1_8 ( .A(new_wire_25), .B(new_wire_451), .C(_1208_), .D(_1206_), .Y(_1209_) );
NOR2X1 NOR2X1_70 ( .A(_788_), .B(_1106_), .Y(_1210_) );
NAND2X1 NAND2X1_81 ( .A(new_wire_218), .B(_1210_), .Y(_1211_) );
INVX1 INVX1_41 ( .A(write_back), .Y(_1212_) );
AND2X2 AND2X2_13 ( .A(_1207_), .B(_1212_), .Y(_1213_) );
NAND2X1 NAND2X1_82 ( .A(new_wire_25), .B(_1213_), .Y(_1214_) );
NOR2X1 NOR2X1_71 ( .A(_1214_), .B(_1211_), .Y(_1215_) );
OR2X2 OR2X2_5 ( .A(_1215_), .B(_1209_), .Y(_1216_) );
NOR2X1 NOR2X1_72 ( .A(_1204_), .B(_1216_), .Y(_1217_) );
OR2X2 OR2X2_6 ( .A(_1194_), .B(_1198_), .Y(_1218_) );
NAND3X1 NAND3X1_49 ( .A(new_wire_22), .B(_1212_), .C(_1218_), .Y(_1219_) );
NAND3X1 NAND3X1_50 ( .A(_1200_), .B(_1219_), .C(_1217_), .Y(_1220_) );
AOI21X1 AOI21X1_39 ( .A(_1189_), .B(new_wire_154), .C(_1220_), .Y(_1221_) );
NAND2X1 NAND2X1_83 ( .A(_1103_), .B(new_wire_403), .Y(_1222_) );
OAI21X1 OAI21X1_72 ( .A(_1089_), .B(new_wire_412), .C(_830__bF_buf2), .Y(_1223_) );
NAND2X1 NAND2X1_84 ( .A(new_wire_395), .B(IRHOLD_6_), .Y(_1224_) );
OAI21X1 OAI21X1_73 ( .A(new_wire_396), .B(new_wire_382), .C(_1224_), .Y(_1225_) );
NAND2X1 NAND2X1_85 ( .A(_830__bF_buf1), .B(_1225_), .Y(_1226_) );
NOR2X1 NOR2X1_73 ( .A(new_wire_453), .B(new_wire_415), .Y(_1227_) );
NAND2X1 NAND2X1_86 ( .A(_1223_), .B(_1227_), .Y(_1228_) );
NOR3X1 NOR3X1_5 ( .A(new_wire_80), .B(_1228_), .C(_1222_), .Y(_1229_) );
NAND3X1 NAND3X1_51 ( .A(_791_), .B(new_wire_253), .C(_801_), .Y(_1230_) );
NOR2X1 NOR2X1_74 ( .A(new_wire_14), .B(_1230_), .Y(_1231_) );
OAI21X1 OAI21X1_74 ( .A(_1207_), .B(_1206_), .C(new_wire_26), .Y(_1232_) );
OAI21X1 OAI21X1_75 ( .A(new_wire_130), .B(_921_), .C(new_wire_189), .Y(_1233_) );
AND2X2 AND2X2_14 ( .A(_1232_), .B(_1233_), .Y(_1234_) );
NOR3X1 NOR3X1_6 ( .A(_1231_), .B(_1234_), .C(_1229_), .Y(_1235_) );
NAND2X1 NAND2X1_87 ( .A(new_wire_338), .B(new_wire_236), .Y(_1236_) );
NOR2X1 NOR2X1_75 ( .A(new_wire_455), .B(new_wire_34), .Y(_1237_) );
NAND2X1 NAND2X1_88 ( .A(new_wire_179), .B(_1237_), .Y(_1238_) );
NAND3X1 NAND3X1_52 ( .A(new_wire_22), .B(write_back), .C(_1218_), .Y(_1239_) );
NOR2X1 NOR2X1_76 ( .A(new_wire_455), .B(new_wire_136), .Y(_1240_) );
OAI21X1 OAI21X1_76 ( .A(new_wire_136), .B(new_wire_339), .C(new_wire_14), .Y(_1241_) );
OAI21X1 OAI21X1_77 ( .A(new_wire_2), .B(_1240_), .C(_1241_), .Y(_1242_) );
NAND3X1 NAND3X1_53 ( .A(_1238_), .B(_1242_), .C(_1239_), .Y(_1243_) );
NAND3X1 NAND3X1_54 ( .A(new_wire_256), .B(new_wire_266), .C(new_wire_247), .Y(_1244_) );
INVX2 INVX2_27 ( .A(_1244_), .Y(_1245_) );
OAI21X1 OAI21X1_78 ( .A(new_wire_138), .B(_803_), .C(new_wire_194), .Y(_1246_) );
OAI21X1 OAI21X1_79 ( .A(new_wire_194), .B(_1245_), .C(_1246_), .Y(_1247_) );
NOR2X1 NOR2X1_77 ( .A(new_wire_227), .B(new_wire_339), .Y(_1248_) );
OAI21X1 OAI21X1_80 ( .A(new_wire_227), .B(new_wire_455), .C(new_wire_182), .Y(_1249_) );
OAI21X1 OAI21X1_81 ( .A(new_wire_182), .B(_1248_), .C(_1249_), .Y(_1250_) );
NOR2X1 NOR2X1_78 ( .A(new_wire_130), .B(new_wire_431), .Y(_1251_) );
OAI21X1 OAI21X1_82 ( .A(new_wire_136), .B(new_wire_427), .C(new_wire_182), .Y(_1252_) );
OAI21X1 OAI21X1_83 ( .A(new_wire_182), .B(new_wire_457), .C(_1252_), .Y(_1253_) );
NAND3X1 NAND3X1_55 ( .A(_1247_), .B(_1250_), .C(_1253_), .Y(_1254_) );
NOR2X1 NOR2X1_79 ( .A(_1254_), .B(_1243_), .Y(_1255_) );
NAND3X1 NAND3X1_56 ( .A(_1255_), .B(_1235_), .C(_1221_), .Y(_1256_) );
NOR2X1 NOR2X1_80 ( .A(_1177_), .B(_1256_), .Y(_1257_) );
NAND3X1 NAND3X1_57 ( .A(_1098_), .B(_1135_), .C(_1257_), .Y(_1438__0_) );
INVX1 INVX1_42 ( .A(_1243_), .Y(_1258_) );
NAND3X1 NAND3X1_58 ( .A(_1250_), .B(_1253_), .C(_1258_), .Y(_1259_) );
NOR2X1 NOR2X1_81 ( .A(_1177_), .B(_1259_), .Y(_1260_) );
NAND2X1 NAND2X1_89 ( .A(new_wire_179), .B(new_wire_457), .Y(_1261_) );
INVX1 INVX1_43 ( .A(IRHOLD_0_), .Y(_1262_) );
AOI21X1 AOI21X1_40 ( .A(new_wire_396), .B(_1262_), .C(new_wire_99), .Y(_1263_) );
OAI21X1 OAI21X1_84 ( .A(new_wire_396), .B(new_wire_374), .C(_1263_), .Y(_1264_) );
OAI21X1 OAI21X1_85 ( .A(new_wire_99), .B(_1082_), .C(_1264_), .Y(_1265_) );
NOR2X1 NOR2X1_82 ( .A(new_wire_459), .B(new_wire_443), .Y(_1266_) );
AND2X2 AND2X2_15 ( .A(_1089_), .B(_830__bF_buf1), .Y(_1267_) );
NAND2X1 NAND2X1_90 ( .A(new_wire_415), .B(new_wire_440), .Y(_1268_) );
NOR2X1 NOR2X1_83 ( .A(new_wire_463), .B(_1268_), .Y(_1269_) );
NAND3X1 NAND3X1_59 ( .A(new_wire_160), .B(_1269_), .C(new_wire_461), .Y(_1270_) );
OAI21X1 OAI21X1_86 ( .A(new_wire_34), .B(new_wire_431), .C(new_wire_179), .Y(_1271_) );
OAI21X1 OAI21X1_87 ( .A(new_wire_179), .B(_1237_), .C(_1271_), .Y(_1272_) );
NAND3X1 NAND3X1_60 ( .A(_1261_), .B(_1272_), .C(_1270_), .Y(_1273_) );
NAND2X1 NAND2X1_91 ( .A(new_wire_407), .B(new_wire_440), .Y(_1274_) );
AND2X2 AND2X2_16 ( .A(_1225_), .B(_830__bF_buf1), .Y(_1275_) );
OAI21X1 OAI21X1_88 ( .A(new_wire_106), .B(new_wire_413), .C(new_wire_467), .Y(_1276_) );
NOR2X1 NOR2X1_84 ( .A(_1276_), .B(new_wire_465), .Y(_1277_) );
NAND2X1 NAND2X1_92 ( .A(new_wire_399), .B(_1181_), .Y(_1278_) );
NOR2X1 NOR2X1_85 ( .A(new_wire_459), .B(_1278_), .Y(_1279_) );
AND2X2 AND2X2_17 ( .A(new_wire_469), .B(_1277_), .Y(_1280_) );
OAI21X1 OAI21X1_89 ( .A(new_wire_135), .B(_806_), .C(new_wire_341), .Y(_1281_) );
NAND2X1 NAND2X1_93 ( .A(new_wire_20), .B(_1281_), .Y(_1282_) );
OAI21X1 OAI21X1_90 ( .A(new_wire_20), .B(_1150_), .C(_1282_), .Y(_1283_) );
AOI21X1 AOI21X1_41 ( .A(_1280_), .B(new_wire_154), .C(_1283_), .Y(_1284_) );
NOR2X1 NOR2X1_86 ( .A(new_wire_227), .B(new_wire_432), .Y(_1285_) );
NAND2X1 NAND2X1_94 ( .A(new_wire_180), .B(_1285_), .Y(_1286_) );
NOR2X1 NOR2X1_87 ( .A(new_wire_445), .B(_1186_), .Y(_1287_) );
AND2X2 AND2X2_18 ( .A(new_wire_471), .B(new_wire_440), .Y(_1288_) );
NAND2X1 NAND2X1_95 ( .A(new_wire_154), .B(_1288_), .Y(_1289_) );
NAND3X1 NAND3X1_61 ( .A(_1286_), .B(_1289_), .C(_1284_), .Y(_1290_) );
NOR2X1 NOR2X1_88 ( .A(new_wire_130), .B(new_wire_438), .Y(_1291_) );
NAND2X1 NAND2X1_96 ( .A(new_wire_453), .B(new_wire_415), .Y(_1292_) );
INVX1 INVX1_44 ( .A(_1292_), .Y(_1293_) );
NAND2X1 NAND2X1_97 ( .A(_1223_), .B(_1293_), .Y(_1294_) );
NOR2X1 NOR2X1_89 ( .A(_1222_), .B(new_wire_476), .Y(_1295_) );
AOI22X1 AOI22X1_16 ( .A(new_wire_176), .B(new_wire_473), .C(new_wire_156), .D(_1295_), .Y(_1296_) );
INVX1 INVX1_45 ( .A(_1160_), .Y(_1297_) );
NOR2X1 NOR2X1_90 ( .A(new_wire_459), .B(_1186_), .Y(_1298_) );
NAND2X1 NAND2X1_98 ( .A(new_wire_467), .B(new_wire_416), .Y(_1299_) );
NOR2X1 NOR2X1_91 ( .A(_1299_), .B(new_wire_465), .Y(_1300_) );
AND2X2 AND2X2_19 ( .A(new_wire_478), .B(new_wire_480), .Y(_1301_) );
AOI22X1 AOI22X1_17 ( .A(new_wire_176), .B(_1297_), .C(new_wire_156), .D(_1301_), .Y(_1302_) );
INVX1 INVX1_46 ( .A(Z), .Y(_1303_) );
NAND2X1 NAND2X1_99 ( .A(new_wire_482), .B(_1303_), .Y(_1304_) );
OAI21X1 OAI21X1_91 ( .A(new_wire_482), .B(C), .C(_1304_), .Y(_1305_) );
INVX2 INVX2_28 ( .A(V), .Y(_1306_) );
NAND2X1 NAND2X1_100 ( .A(new_wire_482), .B(_1306_), .Y(_1307_) );
OAI21X1 OAI21X1_92 ( .A(new_wire_482), .B(N), .C(_1307_), .Y(_1308_) );
MUX2X1 MUX2X1_9 ( .A(_1305_), .B(_1308_), .S(cond_code_2_), .Y(_1309_) );
XNOR2X1 XNOR2X1_1 ( .A(_1309_), .B(cond_code_0_), .Y(_1310_) );
NAND3X1 NAND3X1_62 ( .A(new_wire_26), .B(_1099_), .C(_1310_), .Y(_1311_) );
INVX1 INVX1_47 ( .A(_1230_), .Y(_1312_) );
NAND2X1 NAND2X1_101 ( .A(new_wire_5), .B(_1312_), .Y(_1313_) );
OAI21X1 OAI21X1_93 ( .A(new_wire_15), .B(_1154_), .C(_1313_), .Y(_1314_) );
AOI21X1 AOI21X1_42 ( .A(new_wire_189), .B(new_wire_86), .C(_1314_), .Y(_1315_) );
AND2X2 AND2X2_20 ( .A(_1311_), .B(_1315_), .Y(_1316_) );
NAND3X1 NAND3X1_63 ( .A(_1316_), .B(_1302_), .C(_1296_), .Y(_1317_) );
NOR3X1 NOR3X1_7 ( .A(_1273_), .B(_1290_), .C(_1317_), .Y(_1318_) );
INVX1 INVX1_48 ( .A(new_wire_339), .Y(_1319_) );
NAND2X1 NAND2X1_102 ( .A(new_wire_247), .B(_1319_), .Y(_1320_) );
OR2X2 OR2X2_7 ( .A(_1320_), .B(new_wire_22), .Y(_1321_) );
NAND3X1 NAND3X1_64 ( .A(new_wire_421), .B(new_wire_154), .C(new_wire_471), .Y(_1322_) );
NOR2X1 NOR2X1_92 ( .A(new_wire_32), .B(new_wire_340), .Y(_1323_) );
OAI21X1 OAI21X1_94 ( .A(new_wire_38), .B(new_wire_390), .C(new_wire_2), .Y(_1324_) );
OAI21X1 OAI21X1_95 ( .A(new_wire_2), .B(new_wire_484), .C(_1324_), .Y(_1325_) );
NAND2X1 NAND2X1_103 ( .A(new_wire_190), .B(new_wire_304), .Y(_1326_) );
OAI21X1 OAI21X1_96 ( .A(new_wire_190), .B(_1122_), .C(_1326_), .Y(_1327_) );
AOI21X1 AOI21X1_43 ( .A(new_wire_183), .B(_1248_), .C(_1327_), .Y(_1328_) );
NAND2X1 NAND2X1_104 ( .A(_1325_), .B(_1328_), .Y(_1329_) );
OAI21X1 OAI21X1_97 ( .A(new_wire_445), .B(new_wire_443), .C(_1278_), .Y(_1330_) );
NOR2X1 NOR2X1_93 ( .A(new_wire_80), .B(new_wire_441), .Y(_1331_) );
AOI21X1 AOI21X1_44 ( .A(_1330_), .B(_1331_), .C(_1329_), .Y(_1332_) );
NAND3X1 NAND3X1_65 ( .A(_1321_), .B(_1322_), .C(_1332_), .Y(_1333_) );
INVX1 INVX1_49 ( .A(_1333_), .Y(_1334_) );
NAND3X1 NAND3X1_66 ( .A(_1260_), .B(_1334_), .C(_1318_), .Y(_1438__1_) );
OAI21X1 OAI21X1_98 ( .A(new_wire_228), .B(_811_), .C(new_wire_180), .Y(_1335_) );
NOR2X1 NOR2X1_94 ( .A(new_wire_244), .B(new_wire_242), .Y(_1336_) );
AOI21X1 AOI21X1_45 ( .A(new_wire_253), .B(_841_), .C(_1336_), .Y(_1337_) );
INVX1 INVX1_50 ( .A(new_wire_451), .Y(_1338_) );
NOR2X1 NOR2X1_95 ( .A(new_wire_484), .B(_1338_), .Y(_1339_) );
OAI21X1 OAI21X1_99 ( .A(new_wire_449), .B(_924_), .C(new_wire_253), .Y(_1340_) );
NAND3X1 NAND3X1_67 ( .A(_1340_), .B(_1337_), .C(_1339_), .Y(_1341_) );
NOR2X1 NOR2X1_96 ( .A(_912_), .B(new_wire_207), .Y(_1342_) );
NOR2X1 NOR2X1_97 ( .A(new_wire_177), .B(_1342_), .Y(_1343_) );
OAI21X1 OAI21X1_100 ( .A(new_wire_418), .B(_1310_), .C(_1343_), .Y(_1344_) );
OR2X2 OR2X2_8 ( .A(_1344_), .B(_1341_), .Y(_1345_) );
NOR2X1 NOR2X1_98 ( .A(new_wire_429), .B(_1181_), .Y(_1346_) );
NOR2X1 NOR2X1_99 ( .A(new_wire_76), .B(_1346_), .Y(_1347_) );
OAI21X1 OAI21X1_101 ( .A(_1096_), .B(new_wire_405), .C(_1347_), .Y(_1348_) );
OAI21X1 OAI21X1_102 ( .A(new_wire_421), .B(_1277_), .C(new_wire_478), .Y(_1349_) );
NOR2X1 NOR2X1_100 ( .A(_1292_), .B(new_wire_465), .Y(_1350_) );
AOI22X1 AOI22X1_18 ( .A(new_wire_469), .B(_1277_), .C(new_wire_478), .D(_1350_), .Y(_1351_) );
AOI22X1 AOI22X1_19 ( .A(new_wire_471), .B(new_wire_441), .C(new_wire_478), .D(new_wire_480), .Y(_1352_) );
NAND3X1 NAND3X1_68 ( .A(_1349_), .B(_1351_), .C(_1352_), .Y(_1353_) );
NOR2X1 NOR2X1_101 ( .A(_1348_), .B(_1353_), .Y(_1354_) );
OAI21X1 OAI21X1_103 ( .A(new_wire_101), .B(new_wire_401), .C(new_wire_463), .Y(_1355_) );
NOR2X1 NOR2X1_102 ( .A(new_wire_422), .B(_1355_), .Y(_1356_) );
AOI22X1 AOI22X1_20 ( .A(_1356_), .B(_1103_), .C(new_wire_441), .D(_1184_), .Y(_1357_) );
OAI21X1 OAI21X1_104 ( .A(new_wire_101), .B(new_wire_401), .C(_1083_), .Y(_1358_) );
NOR2X1 NOR2X1_103 ( .A(new_wire_486), .B(new_wire_443), .Y(_1359_) );
AOI21X1 AOI21X1_46 ( .A(new_wire_461), .B(new_wire_465), .C(_1359_), .Y(_1360_) );
OR2X2 OR2X2_9 ( .A(new_wire_413), .B(new_wire_106), .Y(_1361_) );
NOR2X1 NOR2X1_104 ( .A(new_wire_463), .B(_1361_), .Y(_1362_) );
NOR3X1 NOR3X1_8 ( .A(new_wire_422), .B(new_wire_459), .C(new_wire_444), .Y(_1363_) );
AOI22X1 AOI22X1_21 ( .A(new_wire_422), .B(_1330_), .C(_1362_), .D(_1363_), .Y(_1364_) );
NAND3X1 NAND3X1_69 ( .A(_1357_), .B(_1360_), .C(_1364_), .Y(_1365_) );
AOI21X1 AOI21X1_47 ( .A(_1292_), .B(new_wire_407), .C(new_wire_422), .Y(_1366_) );
NAND2X1 NAND2X1_105 ( .A(new_wire_486), .B(new_wire_445), .Y(_1367_) );
NOR2X1 NOR2X1_105 ( .A(new_wire_423), .B(_1278_), .Y(_1368_) );
AOI22X1 AOI22X1_22 ( .A(new_wire_469), .B(_1366_), .C(_1367_), .D(_1368_), .Y(_1369_) );
OAI21X1 OAI21X1_105 ( .A(_1089_), .B(_1225_), .C(new_wire_165), .Y(_1370_) );
NAND3X1 NAND3X1_70 ( .A(_1095_), .B(_1370_), .C(new_wire_479), .Y(_1371_) );
AOI22X1 AOI22X1_23 ( .A(new_wire_469), .B(new_wire_480), .C(new_wire_423), .D(new_wire_471), .Y(_1372_) );
NAND3X1 NAND3X1_71 ( .A(_1371_), .B(_1369_), .C(_1372_), .Y(_1373_) );
NOR2X1 NOR2X1_106 ( .A(_1373_), .B(_1365_), .Y(_1374_) );
AOI22X1 AOI22X1_24 ( .A(_1335_), .B(_1345_), .C(_1354_), .D(_1374_), .Y(_1375_) );
INVX1 INVX1_51 ( .A(new_wire_449), .Y(_1376_) );
OAI21X1 OAI21X1_106 ( .A(new_wire_136), .B(_1376_), .C(new_wire_183), .Y(_1377_) );
OAI21X1 OAI21X1_107 ( .A(new_wire_183), .B(_1240_), .C(_1377_), .Y(_1378_) );
INVX1 INVX1_52 ( .A(_1378_), .Y(_1379_) );
OAI21X1 OAI21X1_108 ( .A(new_wire_138), .B(new_wire_436), .C(new_wire_15), .Y(_1380_) );
OAI21X1 OAI21X1_109 ( .A(new_wire_15), .B(_1245_), .C(_1380_), .Y(_1381_) );
OAI21X1 OAI21X1_110 ( .A(new_wire_37), .B(new_wire_436), .C(new_wire_21), .Y(_1382_) );
OAI21X1 OAI21X1_111 ( .A(new_wire_21), .B(_1202_), .C(_1382_), .Y(_1383_) );
NAND2X1 NAND2X1_106 ( .A(_1383_), .B(_1381_), .Y(_1384_) );
NOR2X1 NOR2X1_107 ( .A(_1384_), .B(_1379_), .Y(_1385_) );
AND2X2 AND2X2_21 ( .A(_1375_), .B(_1385_), .Y(_1386_) );
OR2X2 OR2X2_10 ( .A(_1290_), .B(_1273_), .Y(_1387_) );
INVX2 INVX2_29 ( .A(new_wire_486), .Y(_1388_) );
NAND2X1 NAND2X1_107 ( .A(_1081_), .B(new_wire_488), .Y(_1389_) );
OAI21X1 OAI21X1_112 ( .A(_1223_), .B(new_wire_405), .C(new_wire_490), .Y(_1390_) );
NAND2X1 NAND2X1_108 ( .A(new_wire_156), .B(_1390_), .Y(_1391_) );
NOR2X1 NOR2X1_108 ( .A(new_wire_39), .B(_1376_), .Y(_1392_) );
NAND2X1 NAND2X1_109 ( .A(new_wire_180), .B(_1392_), .Y(_1393_) );
INVX1 INVX1_53 ( .A(_1197_), .Y(_1394_) );
OAI21X1 OAI21X1_113 ( .A(_1213_), .B(_1211_), .C(new_wire_23), .Y(_1395_) );
OAI21X1 OAI21X1_114 ( .A(new_wire_23), .B(_1394_), .C(_1395_), .Y(_1396_) );
NAND3X1 NAND3X1_72 ( .A(_1393_), .B(_1396_), .C(_1391_), .Y(_1397_) );
NAND3X1 NAND3X1_73 ( .A(_1247_), .B(_1253_), .C(_1169_), .Y(_1398_) );
NOR2X1 NOR2X1_109 ( .A(_1398_), .B(_1105_), .Y(_1399_) );
NAND3X1 NAND3X1_74 ( .A(_1316_), .B(_1159_), .C(_1399_), .Y(_1400_) );
NOR2X1 NOR2X1_110 ( .A(_1397_), .B(_1400_), .Y(_1401_) );
NAND3X1 NAND3X1_75 ( .A(_1221_), .B(_1235_), .C(_1401_), .Y(_1402_) );
NOR2X1 NOR2X1_111 ( .A(_1387_), .B(_1402_), .Y(_1403_) );
NAND2X1 NAND2X1_110 ( .A(_1386_), .B(_1403_), .Y(_1438__2_) );
INVX1 INVX1_54 ( .A(_1127_), .Y(_1404_) );
NAND3X1 NAND3X1_76 ( .A(new_wire_155), .B(new_wire_480), .C(new_wire_470), .Y(_1405_) );
OAI21X1 OAI21X1_115 ( .A(new_wire_23), .B(_1404_), .C(_1405_), .Y(_1406_) );
OAI21X1 OAI21X1_116 ( .A(new_wire_34), .B(new_wire_425), .C(new_wire_183), .Y(_1407_) );
OAI21X1 OAI21X1_117 ( .A(new_wire_35), .B(new_wire_242), .C(new_wire_2), .Y(_1408_) );
AOI21X1 AOI21X1_48 ( .A(_1407_), .B(_1408_), .C(_1406_), .Y(_1409_) );
INVX1 INVX1_55 ( .A(_1409_), .Y(_1410_) );
AOI22X1 AOI22X1_25 ( .A(new_wire_180), .B(_1111_), .C(_1331_), .D(_1346_), .Y(_1411_) );
OAI21X1 OAI21X1_118 ( .A(_923_), .B(new_wire_137), .C(new_wire_184), .Y(_1412_) );
OAI21X1 OAI21X1_119 ( .A(new_wire_181), .B(_1144_), .C(_1412_), .Y(_1413_) );
NAND2X1 NAND2X1_111 ( .A(_1413_), .B(_1411_), .Y(_1414_) );
NAND2X1 NAND2X1_112 ( .A(new_wire_213), .B(_924_), .Y(_1415_) );
NOR2X1 NOR2X1_112 ( .A(_923_), .B(new_wire_35), .Y(_1416_) );
OAI21X1 OAI21X1_120 ( .A(new_wire_130), .B(new_wire_427), .C(new_wire_3), .Y(_1417_) );
OAI21X1 OAI21X1_121 ( .A(new_wire_3), .B(_1416_), .C(_1417_), .Y(_1418_) );
OAI21X1 OAI21X1_122 ( .A(new_wire_3), .B(_1415_), .C(_1418_), .Y(_1419_) );
NOR2X1 NOR2X1_113 ( .A(_1419_), .B(_1414_), .Y(_1420_) );
OAI21X1 OAI21X1_123 ( .A(new_wire_76), .B(_1369_), .C(_1420_), .Y(_1421_) );
NOR2X1 NOR2X1_114 ( .A(_1421_), .B(_1410_), .Y(_1422_) );
NAND2X1 NAND2X1_113 ( .A(_1098_), .B(_1135_), .Y(_1423_) );
NOR3X1 NOR3X1_9 ( .A(_1333_), .B(_1397_), .C(_1423_), .Y(_1424_) );
NAND3X1 NAND3X1_77 ( .A(_1422_), .B(_1424_), .C(_1318_), .Y(_1425_) );
NAND3X1 NAND3X1_78 ( .A(_1385_), .B(_1375_), .C(_1257_), .Y(_1426_) );
OAI21X1 OAI21X1_124 ( .A(_1341_), .B(_1344_), .C(_1335_), .Y(_1427_) );
NAND2X1 NAND2X1_114 ( .A(_1354_), .B(_1374_), .Y(_1428_) );
NAND2X1 NAND2X1_115 ( .A(_1427_), .B(_1428_), .Y(_1429_) );
NAND2X1 NAND2X1_116 ( .A(new_wire_441), .B(new_wire_472), .Y(_1430_) );
OAI21X1 OAI21X1_125 ( .A(new_wire_76), .B(_1430_), .C(_1286_), .Y(_1431_) );
NAND2X1 NAND2X1_117 ( .A(_1173_), .B(_1253_), .Y(_1432_) );
NAND2X1 NAND2X1_118 ( .A(_1247_), .B(_1129_), .Y(_1433_) );
NOR2X1 NOR2X1_115 ( .A(_1433_), .B(_1432_), .Y(_1434_) );
OR2X2 OR2X2_11 ( .A(_1125_), .B(_1121_), .Y(_1435_) );
NOR2X1 NOR2X1_116 ( .A(_1327_), .B(_1435_), .Y(_1436_) );
NOR2X1 NOR2X1_117 ( .A(_1384_), .B(_1166_), .Y(_1437_) );
NAND3X1 NAND3X1_79 ( .A(_1434_), .B(_1437_), .C(_1436_), .Y(_41_) );
NOR3X1 NOR3X1_10 ( .A(_1148_), .B(_1431_), .C(_41_), .Y(_42_) );
INVX2 INVX2_30 ( .A(new_wire_473), .Y(_43_) );
NAND2X1 NAND2X1_119 ( .A(_1350_), .B(new_wire_479), .Y(_44_) );
OAI22X1 OAI22X1_9 ( .A(new_wire_23), .B(new_wire_492), .C(new_wire_77), .D(_44_), .Y(_45_) );
NAND2X1 NAND2X1_120 ( .A(new_wire_481), .B(new_wire_479), .Y(_46_) );
OAI22X1 OAI22X1_10 ( .A(new_wire_24), .B(_1160_), .C(new_wire_77), .D(_46_), .Y(_47_) );
NOR3X1 NOR3X1_11 ( .A(_1273_), .B(_45_), .C(_47_), .Y(_48_) );
AND2X2 AND2X2_22 ( .A(_1221_), .B(_1409_), .Y(_49_) );
NAND3X1 NAND3X1_80 ( .A(_42_), .B(_48_), .C(_49_), .Y(_50_) );
NOR2X1 NOR2X1_118 ( .A(_50_), .B(_1429_), .Y(_51_) );
OAI21X1 OAI21X1_126 ( .A(_1425_), .B(_1426_), .C(_51_), .Y(_1438__3_) );
INVX1 INVX1_56 ( .A(_1234_), .Y(_52_) );
NAND3X1 NAND3X1_81 ( .A(_1117_), .B(_1152_), .C(_52_), .Y(_53_) );
AND2X2 AND2X2_23 ( .A(_1242_), .B(_1381_), .Y(_54_) );
NAND3X1 NAND3X1_82 ( .A(_1378_), .B(_54_), .C(_1434_), .Y(_55_) );
OR2X2 OR2X2_12 ( .A(_55_), .B(_53_), .Y(_56_) );
NOR2X1 NOR2X1_119 ( .A(_45_), .B(_56_), .Y(_57_) );
OAI21X1 OAI21X1_127 ( .A(new_wire_24), .B(_1320_), .C(_1322_), .Y(_58_) );
NOR2X1 NOR2X1_120 ( .A(_1414_), .B(_58_), .Y(_59_) );
NAND3X1 NAND3X1_83 ( .A(_1261_), .B(_1270_), .C(_1284_), .Y(_60_) );
NOR2X1 NOR2X1_121 ( .A(_1406_), .B(_60_), .Y(_61_) );
NAND3X1 NAND3X1_84 ( .A(_57_), .B(_59_), .C(_61_), .Y(_1438__4_) );
AND2X2 AND2X2_24 ( .A(_1239_), .B(_1238_), .Y(_62_) );
INVX1 INVX1_57 ( .A(_1325_), .Y(_63_) );
NOR2X1 NOR2X1_122 ( .A(_1314_), .B(_63_), .Y(_64_) );
INVX1 INVX1_58 ( .A(_1272_), .Y(_65_) );
NOR2X1 NOR2X1_123 ( .A(_1164_), .B(_65_), .Y(_66_) );
NOR2X1 NOR2X1_124 ( .A(_1121_), .B(_1113_), .Y(_67_) );
NOR2X1 NOR2X1_125 ( .A(_1204_), .B(_1157_), .Y(_68_) );
AND2X2 AND2X2_25 ( .A(_68_), .B(_67_), .Y(_69_) );
NAND3X1 NAND3X1_85 ( .A(_64_), .B(_66_), .C(_69_), .Y(_70_) );
INVX1 INVX1_59 ( .A(_1418_), .Y(_71_) );
AOI21X1 AOI21X1_49 ( .A(_1407_), .B(_1408_), .C(_71_), .Y(_72_) );
NAND3X1 NAND3X1_86 ( .A(_1142_), .B(_1383_), .C(_72_), .Y(_73_) );
NOR2X1 NOR2X1_126 ( .A(_73_), .B(_70_), .Y(_74_) );
NAND3X1 NAND3X1_87 ( .A(_62_), .B(_1411_), .C(_74_), .Y(_75_) );
NOR2X1 NOR2X1_127 ( .A(_1231_), .B(_1229_), .Y(_76_) );
NAND3X1 NAND3X1_88 ( .A(_1098_), .B(_1302_), .C(_76_), .Y(_77_) );
NOR2X1 NOR2X1_128 ( .A(_77_), .B(_75_), .Y(_78_) );
NAND3X1 NAND3X1_89 ( .A(_1391_), .B(_1393_), .C(_78_), .Y(_1438__5_) );
INVX1 INVX1_60 ( .A(C), .Y(_79_) );
OAI21X1 OAI21X1_128 ( .A(new_wire_450), .B(_1210_), .C(new_wire_253), .Y(_80_) );
OAI21X1 OAI21X1_129 ( .A(_803_), .B(new_wire_225), .C(_80_), .Y(_81_) );
OR2X2 OR2X2_13 ( .A(new_wire_451), .B(load_only), .Y(_82_) );
NOR2X1 NOR2X1_129 ( .A(shift), .B(_82_), .Y(_83_) );
AOI21X1 AOI21X1_50 ( .A(rotate), .B(new_wire_494), .C(_83_), .Y(_84_) );
INVX1 INVX1_61 ( .A(rotate), .Y(_85_) );
INVX2 INVX2_31 ( .A(compare), .Y(_86_) );
INVX2 INVX2_32 ( .A(shift), .Y(_87_) );
INVX1 INVX1_62 ( .A(_80_), .Y(_88_) );
NAND3X1 NAND3X1_90 ( .A(inc), .B(_87_), .C(_88_), .Y(_89_) );
OAI21X1 OAI21X1_130 ( .A(new_wire_496), .B(new_wire_451), .C(_89_), .Y(_90_) );
INVX1 INVX1_63 ( .A(_1206_), .Y(_91_) );
OAI21X1 OAI21X1_131 ( .A(new_wire_223), .B(new_wire_455), .C(new_wire_207), .Y(_92_) );
OAI21X1 OAI21X1_132 ( .A(_91_), .B(_92_), .C(new_wire_335), .Y(_93_) );
OAI21X1 OAI21X1_133 ( .A(new_wire_30), .B(new_wire_437), .C(_1154_), .Y(_94_) );
OAI21X1 OAI21X1_134 ( .A(new_wire_30), .B(new_wire_438), .C(_1230_), .Y(_95_) );
OR2X2 OR2X2_14 ( .A(_94_), .B(_95_), .Y(_96_) );
INVX1 INVX1_64 ( .A(new_wire_457), .Y(_97_) );
OAI21X1 OAI21X1_135 ( .A(new_wire_32), .B(new_wire_242), .C(_1143_), .Y(_98_) );
INVX1 INVX1_65 ( .A(_98_), .Y(_99_) );
NAND3X1 NAND3X1_91 ( .A(_1320_), .B(_97_), .C(_99_), .Y(_100_) );
NOR2X1 NOR2X1_130 ( .A(_100_), .B(_96_), .Y(_101_) );
NAND2X1 NAND2X1_121 ( .A(_93_), .B(_101_), .Y(_102_) );
AOI21X1 AOI21X1_51 ( .A(_85_), .B(_90_), .C(_102_), .Y(_103_) );
OAI21X1 OAI21X1_136 ( .A(_79_), .B(_84_), .C(_103_), .Y(CI) );
INVX2 INVX2_33 ( .A(new_wire_374), .Y(_104_) );
NOR2X1 NOR2X1_131 ( .A(new_wire_473), .B(_88_), .Y(_105_) );
AOI21X1 AOI21X1_52 ( .A(_841_), .B(new_wire_214), .C(_1170_), .Y(_106_) );
NOR2X1 NOR2X1_132 ( .A(new_wire_87), .B(_1245_), .Y(_107_) );
NAND2X1 NAND2X1_122 ( .A(_107_), .B(new_wire_498), .Y(_108_) );
NOR2X1 NOR2X1_133 ( .A(_840_), .B(_1195_), .Y(_109_) );
OAI21X1 OAI21X1_137 ( .A(new_wire_305), .B(_109_), .C(new_wire_216), .Y(_110_) );
NOR2X1 NOR2X1_134 ( .A(new_wire_392), .B(new_wire_457), .Y(_111_) );
NAND2X1 NAND2X1_123 ( .A(_110_), .B(_111_), .Y(_112_) );
NOR2X1 NOR2X1_135 ( .A(_108_), .B(_112_), .Y(_113_) );
INVX2 INVX2_34 ( .A(new_wire_484), .Y(_114_) );
NAND3X1 NAND3X1_92 ( .A(new_wire_500), .B(_99_), .C(new_wire_418), .Y(_115_) );
NOR2X1 NOR2X1_136 ( .A(_96_), .B(_115_), .Y(_116_) );
NAND3X1 NAND3X1_93 ( .A(_105_), .B(_113_), .C(_116_), .Y(_117_) );
OAI22X1 OAI22X1_11 ( .A(new_wire_333), .B(new_wire_418), .C(_104_), .D(new_wire_502), .Y(BI_0_) );
INVX2 INVX2_35 ( .A(new_wire_372), .Y(_118_) );
OAI22X1 OAI22X1_12 ( .A(new_wire_349), .B(new_wire_419), .C(_118_), .D(new_wire_502), .Y(BI_1_) );
OAI22X1 OAI22X1_13 ( .A(new_wire_360), .B(new_wire_419), .C(new_wire_366), .D(new_wire_502), .Y(BI_2_) );
OAI22X1 OAI22X1_14 ( .A(new_wire_354), .B(new_wire_419), .C(_1179_), .D(new_wire_502), .Y(BI_3_) );
OAI22X1 OAI22X1_15 ( .A(new_wire_318), .B(new_wire_419), .C(new_wire_378), .D(new_wire_503), .Y(BI_4_) );
INVX1 INVX1_66 ( .A(new_wire_293), .Y(_119_) );
OAI22X1 OAI22X1_16 ( .A(new_wire_307), .B(new_wire_420), .C(_119_), .D(new_wire_503), .Y(BI_5_) );
OAI22X1 OAI22X1_17 ( .A(new_wire_328), .B(new_wire_420), .C(new_wire_382), .D(new_wire_503), .Y(BI_6_) );
OAI22X1 OAI22X1_18 ( .A(new_wire_323), .B(new_wire_420), .C(new_wire_386), .D(new_wire_503), .Y(BI_7_) );
NOR2X1 NOR2X1_137 ( .A(_1006_), .B(new_wire_203), .Y(_120_) );
OAI21X1 OAI21X1_138 ( .A(new_wire_225), .B(new_wire_438), .C(new_wire_498), .Y(_121_) );
OR2X2 OR2X2_15 ( .A(_121_), .B(_94_), .Y(_122_) );
OAI21X1 OAI21X1_139 ( .A(_98_), .B(_122_), .C(new_wire_330), .Y(_123_) );
OAI21X1 OAI21X1_140 ( .A(new_wire_32), .B(new_wire_456), .C(new_wire_420), .Y(_124_) );
INVX4 INVX4_4 ( .A(_124_), .Y(_125_) );
OAI21X1 OAI21X1_141 ( .A(_104_), .B(new_wire_508), .C(_123_), .Y(_126_) );
NOR2X1 NOR2X1_138 ( .A(_120_), .B(_126_), .Y(_127_) );
INVX1 INVX1_67 ( .A(src_reg_1_), .Y(_128_) );
OAI21X1 OAI21X1_142 ( .A(new_wire_230), .B(new_wire_340), .C(_1110_), .Y(_129_) );
OAI22X1 OAI22X1_19 ( .A(new_wire_131), .B(new_wire_456), .C(new_wire_223), .D(new_wire_432), .Y(_130_) );
NOR3X1 NOR3X1_12 ( .A(new_wire_197), .B(_129_), .C(_130_), .Y(_131_) );
OAI22X1 OAI22X1_20 ( .A(new_wire_225), .B(new_wire_426), .C(new_wire_132), .D(new_wire_439), .Y(_132_) );
OAI21X1 OAI21X1_143 ( .A(new_wire_32), .B(new_wire_426), .C(_1160_), .Y(_133_) );
NOR2X1 NOR2X1_139 ( .A(new_wire_510), .B(_133_), .Y(_134_) );
OAI21X1 OAI21X1_144 ( .A(new_wire_131), .B(new_wire_432), .C(new_wire_341), .Y(_135_) );
NAND2X1 NAND2X1_124 ( .A(new_wire_247), .B(_1137_), .Y(_136_) );
OAI21X1 OAI21X1_145 ( .A(new_wire_33), .B(new_wire_340), .C(_136_), .Y(_137_) );
NAND3X1 NAND3X1_94 ( .A(_1201_), .B(_1244_), .C(_1230_), .Y(_138_) );
NOR3X1 NOR3X1_13 ( .A(_137_), .B(_135_), .C(_138_), .Y(_139_) );
NAND3X1 NAND3X1_95 ( .A(_131_), .B(_139_), .C(_134_), .Y(_140_) );
INVX1 INVX1_68 ( .A(dst_reg_1_), .Y(_141_) );
NOR2X1 NOR2X1_140 ( .A(_129_), .B(_130_), .Y(_142_) );
OAI21X1 OAI21X1_146 ( .A(_141_), .B(new_wire_122), .C(_142_), .Y(_143_) );
INVX1 INVX1_69 ( .A(_143_), .Y(_144_) );
OAI21X1 OAI21X1_147 ( .A(_128_), .B(_140_), .C(_144_), .Y(_145_) );
INVX4 INVX4_5 ( .A(new_wire_512), .Y(_146_) );
INVX1 INVX1_70 ( .A(AXYS_1__0_), .Y(_147_) );
OR2X2 OR2X2_16 ( .A(_140_), .B(src_reg_0_), .Y(_148_) );
OAI21X1 OAI21X1_148 ( .A(new_wire_224), .B(_811_), .C(_142_), .Y(_149_) );
OAI21X1 OAI21X1_149 ( .A(_129_), .B(_130_), .C(index_y), .Y(_150_) );
NAND2X1 NAND2X1_125 ( .A(dst_reg_0_), .B(new_wire_197), .Y(_151_) );
NAND3X1 NAND3X1_96 ( .A(_150_), .B(_151_), .C(_149_), .Y(_152_) );
NAND3X1 NAND3X1_97 ( .A(_147_), .B(new_wire_124), .C(_148__bF_buf2), .Y(_153_) );
INVX1 INVX1_71 ( .A(AXYS_0__0_), .Y(_154_) );
OAI21X1 OAI21X1_150 ( .A(src_reg_0_), .B(_140_), .C(_152__bF_buf1), .Y(_155_) );
NAND2X1 NAND2X1_126 ( .A(_154_), .B(_155__bF_buf1), .Y(_156_) );
NAND3X1 NAND3X1_98 ( .A(new_wire_515), .B(_156_), .C(_153_), .Y(_157_) );
INVX1 INVX1_72 ( .A(AXYS_3__0_), .Y(_158_) );
NAND3X1 NAND3X1_99 ( .A(_158_), .B(new_wire_124), .C(_148__bF_buf2), .Y(_159_) );
INVX1 INVX1_73 ( .A(AXYS_2__0_), .Y(_160_) );
NAND2X1 NAND2X1_127 ( .A(_160_), .B(new_wire_108), .Y(_161_) );
NAND3X1 NAND3X1_100 ( .A(new_wire_512), .B(_161_), .C(_159_), .Y(_162_) );
AND2X2 AND2X2_26 ( .A(_157_), .B(_162_), .Y(_163_) );
NOR2X1 NOR2X1_141 ( .A(new_wire_392), .B(_1123_), .Y(_164_) );
OAI21X1 OAI21X1_151 ( .A(new_wire_343), .B(_1319_), .C(new_wire_254), .Y(_165_) );
OAI21X1 OAI21X1_152 ( .A(new_wire_248), .B(new_wire_254), .C(new_wire_306), .Y(_166_) );
AND2X2 AND2X2_27 ( .A(_165_), .B(_166_), .Y(_167_) );
NAND3X1 NAND3X1_101 ( .A(_82_), .B(_164_), .C(_167_), .Y(_168_) );
INVX1 INVX1_74 ( .A(_1392_), .Y(_169_) );
NOR2X1 NOR2X1_142 ( .A(_1245_), .B(new_wire_458), .Y(_170_) );
NAND3X1 NAND3X1_102 ( .A(_169_), .B(_170_), .C(_142_), .Y(_171_) );
NOR2X1 NOR2X1_143 ( .A(_171_), .B(_168_), .Y(_172_) );
OAI21X1 OAI21X1_153 ( .A(new_wire_518), .B(_163_), .C(_127_), .Y(AI_0_) );
OR2X2 OR2X2_17 ( .A(_122_), .B(_98_), .Y(_173_) );
OAI22X1 OAI22X1_21 ( .A(_994_), .B(new_wire_203), .C(_118_), .D(new_wire_508), .Y(_174_) );
AOI21X1 AOI21X1_53 ( .A(new_wire_520), .B(new_wire_345), .C(_174_), .Y(_175_) );
INVX1 INVX1_75 ( .A(AXYS_1__1_), .Y(_176_) );
NAND3X1 NAND3X1_103 ( .A(_176_), .B(_152__bF_buf1), .C(_148__bF_buf0), .Y(_177_) );
INVX1 INVX1_76 ( .A(AXYS_0__1_), .Y(_178_) );
NAND2X1 NAND2X1_128 ( .A(_178_), .B(_155__bF_buf0), .Y(_179_) );
NAND3X1 NAND3X1_104 ( .A(new_wire_515), .B(_179_), .C(_177_), .Y(_180_) );
INVX1 INVX1_77 ( .A(AXYS_3__1_), .Y(_181_) );
NAND3X1 NAND3X1_105 ( .A(_181_), .B(new_wire_124), .C(_148__bF_buf0), .Y(_182_) );
INVX1 INVX1_78 ( .A(AXYS_2__1_), .Y(_183_) );
NAND2X1 NAND2X1_129 ( .A(_183_), .B(new_wire_108), .Y(_184_) );
NAND3X1 NAND3X1_106 ( .A(new_wire_512), .B(_184_), .C(_182_), .Y(_185_) );
AND2X2 AND2X2_28 ( .A(_180_), .B(_185_), .Y(_186_) );
OAI21X1 OAI21X1_154 ( .A(new_wire_518), .B(_186_), .C(_175_), .Y(AI_1_) );
OAI22X1 OAI22X1_22 ( .A(_981_), .B(new_wire_203), .C(new_wire_366), .D(new_wire_508), .Y(_187_) );
AOI21X1 AOI21X1_54 ( .A(new_wire_520), .B(new_wire_357), .C(_187_), .Y(_188_) );
INVX1 INVX1_79 ( .A(AXYS_1__2_), .Y(_189_) );
NAND3X1 NAND3X1_107 ( .A(_189_), .B(new_wire_126), .C(new_wire_201), .Y(_190_) );
INVX1 INVX1_80 ( .A(AXYS_0__2_), .Y(_191_) );
NAND2X1 NAND2X1_130 ( .A(_191_), .B(new_wire_110), .Y(_192_) );
NAND3X1 NAND3X1_108 ( .A(new_wire_515), .B(_192_), .C(_190_), .Y(_193_) );
INVX1 INVX1_81 ( .A(AXYS_3__2_), .Y(_194_) );
NAND3X1 NAND3X1_109 ( .A(_194_), .B(new_wire_126), .C(new_wire_201), .Y(_195_) );
INVX1 INVX1_82 ( .A(AXYS_2__2_), .Y(_196_) );
NAND2X1 NAND2X1_131 ( .A(_196_), .B(new_wire_110), .Y(_197_) );
NAND3X1 NAND3X1_110 ( .A(new_wire_512), .B(_197_), .C(_195_), .Y(_198_) );
AND2X2 AND2X2_29 ( .A(_193_), .B(_198_), .Y(_199_) );
OAI21X1 OAI21X1_155 ( .A(new_wire_518), .B(_199_), .C(_188_), .Y(AI_2_) );
OAI22X1 OAI22X1_23 ( .A(_970_), .B(new_wire_203), .C(_1179_), .D(new_wire_508), .Y(_200_) );
AOI21X1 AOI21X1_55 ( .A(new_wire_520), .B(new_wire_352), .C(_200_), .Y(_201_) );
INVX1 INVX1_83 ( .A(AXYS_1__3_), .Y(_202_) );
NAND3X1 NAND3X1_111 ( .A(_202_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_203_) );
INVX1 INVX1_84 ( .A(AXYS_0__3_), .Y(_204_) );
NAND2X1 NAND2X1_132 ( .A(_204_), .B(new_wire_108), .Y(_205_) );
NAND3X1 NAND3X1_112 ( .A(new_wire_515), .B(_205_), .C(_203_), .Y(_206_) );
INVX1 INVX1_85 ( .A(AXYS_3__3_), .Y(_207_) );
NAND3X1 NAND3X1_113 ( .A(_207_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_208_) );
INVX1 INVX1_86 ( .A(AXYS_2__3_), .Y(_209_) );
NAND2X1 NAND2X1_133 ( .A(_209_), .B(_155__bF_buf0), .Y(_210_) );
NAND3X1 NAND3X1_114 ( .A(new_wire_513), .B(_210_), .C(_208_), .Y(_211_) );
AND2X2 AND2X2_30 ( .A(_206_), .B(_211_), .Y(_212_) );
OAI21X1 OAI21X1_156 ( .A(new_wire_518), .B(_212_), .C(_201_), .Y(AI_3_) );
OAI22X1 OAI22X1_24 ( .A(_1020_), .B(new_wire_204), .C(new_wire_378), .D(new_wire_509), .Y(_213_) );
AOI21X1 AOI21X1_56 ( .A(new_wire_520), .B(new_wire_312), .C(_213_), .Y(_214_) );
INVX1 INVX1_87 ( .A(AXYS_1__4_), .Y(_215_) );
NAND3X1 NAND3X1_115 ( .A(_215_), .B(_152__bF_buf1), .C(_148__bF_buf0), .Y(_216_) );
INVX1 INVX1_88 ( .A(AXYS_0__4_), .Y(_217_) );
NAND2X1 NAND2X1_134 ( .A(_217_), .B(_155__bF_buf0), .Y(_218_) );
NAND3X1 NAND3X1_116 ( .A(new_wire_516), .B(_218_), .C(_216_), .Y(_219_) );
INVX1 INVX1_89 ( .A(AXYS_3__4_), .Y(_220_) );
NAND3X1 NAND3X1_117 ( .A(_220_), .B(_152__bF_buf1), .C(_148__bF_buf0), .Y(_221_) );
INVX1 INVX1_90 ( .A(AXYS_2__4_), .Y(_222_) );
NAND2X1 NAND2X1_135 ( .A(_222_), .B(new_wire_108), .Y(_223_) );
NAND3X1 NAND3X1_118 ( .A(new_wire_513), .B(_223_), .C(_221_), .Y(_224_) );
AND2X2 AND2X2_31 ( .A(_219_), .B(_224_), .Y(_225_) );
OAI21X1 OAI21X1_157 ( .A(new_wire_519), .B(_225_), .C(_214_), .Y(AI_4_) );
INVX1 INVX1_91 ( .A(ABH_5_), .Y(_226_) );
OAI22X1 OAI22X1_25 ( .A(_226_), .B(new_wire_205), .C(_119_), .D(new_wire_509), .Y(_227_) );
AOI21X1 AOI21X1_57 ( .A(new_wire_521), .B(new_wire_295), .C(_227_), .Y(_228_) );
INVX1 INVX1_92 ( .A(AXYS_1__5_), .Y(_229_) );
NAND3X1 NAND3X1_119 ( .A(_229_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_230_) );
INVX1 INVX1_93 ( .A(AXYS_0__5_), .Y(_231_) );
NAND2X1 NAND2X1_136 ( .A(_231_), .B(_155__bF_buf1), .Y(_232_) );
NAND3X1 NAND3X1_120 ( .A(new_wire_516), .B(_232_), .C(_230_), .Y(_233_) );
INVX1 INVX1_94 ( .A(AXYS_3__5_), .Y(_234_) );
NAND3X1 NAND3X1_121 ( .A(_234_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_235_) );
INVX1 INVX1_95 ( .A(AXYS_2__5_), .Y(_236_) );
NAND2X1 NAND2X1_137 ( .A(_236_), .B(new_wire_109), .Y(_237_) );
NAND3X1 NAND3X1_122 ( .A(new_wire_513), .B(_237_), .C(_235_), .Y(_238_) );
AND2X2 AND2X2_32 ( .A(_233_), .B(_238_), .Y(_239_) );
OAI21X1 OAI21X1_158 ( .A(new_wire_519), .B(_239_), .C(_228_), .Y(AI_5_) );
OAI22X1 OAI22X1_26 ( .A(_1049_), .B(new_wire_205), .C(new_wire_382), .D(new_wire_509), .Y(_240_) );
AOI21X1 AOI21X1_58 ( .A(new_wire_521), .B(new_wire_325), .C(_240_), .Y(_241_) );
INVX1 INVX1_96 ( .A(AXYS_1__6_), .Y(_242_) );
NAND3X1 NAND3X1_123 ( .A(_242_), .B(new_wire_124), .C(_148__bF_buf2), .Y(_243_) );
INVX1 INVX1_97 ( .A(AXYS_0__6_), .Y(_244_) );
NAND2X1 NAND2X1_138 ( .A(_244_), .B(_155__bF_buf1), .Y(_245_) );
NAND3X1 NAND3X1_124 ( .A(new_wire_516), .B(_245_), .C(_243_), .Y(_246_) );
INVX1 INVX1_98 ( .A(AXYS_3__6_), .Y(_247_) );
NAND3X1 NAND3X1_125 ( .A(_247_), .B(new_wire_125), .C(_148__bF_buf2), .Y(_248_) );
INVX1 INVX1_99 ( .A(AXYS_2__6_), .Y(_249_) );
NAND2X1 NAND2X1_139 ( .A(_249_), .B(_155__bF_buf1), .Y(_250_) );
NAND3X1 NAND3X1_126 ( .A(new_wire_513), .B(_250_), .C(_248_), .Y(_251_) );
AND2X2 AND2X2_33 ( .A(_246_), .B(_251_), .Y(_252_) );
OAI21X1 OAI21X1_159 ( .A(new_wire_519), .B(_252_), .C(_241_), .Y(AI_6_) );
OAI22X1 OAI22X1_27 ( .A(_1061_), .B(new_wire_205), .C(new_wire_386), .D(new_wire_509), .Y(_253_) );
AOI21X1 AOI21X1_59 ( .A(new_wire_521), .B(new_wire_320), .C(_253_), .Y(_254_) );
INVX1 INVX1_100 ( .A(AXYS_1__7_), .Y(_255_) );
NAND3X1 NAND3X1_127 ( .A(_255_), .B(new_wire_126), .C(new_wire_201), .Y(_256_) );
INVX1 INVX1_101 ( .A(AXYS_0__7_), .Y(_257_) );
NAND2X1 NAND2X1_140 ( .A(_257_), .B(new_wire_110), .Y(_258_) );
NAND3X1 NAND3X1_128 ( .A(new_wire_516), .B(_258_), .C(_256_), .Y(_259_) );
INVX1 INVX1_102 ( .A(AXYS_3__7_), .Y(_260_) );
NAND3X1 NAND3X1_129 ( .A(_260_), .B(new_wire_126), .C(new_wire_201), .Y(_261_) );
INVX1 INVX1_103 ( .A(AXYS_2__7_), .Y(_262_) );
NAND2X1 NAND2X1_141 ( .A(_262_), .B(new_wire_110), .Y(_263_) );
NAND3X1 NAND3X1_130 ( .A(new_wire_514), .B(_263_), .C(_261_), .Y(_264_) );
AND2X2 AND2X2_34 ( .A(_259_), .B(_264_), .Y(_265_) );
OAI21X1 OAI21X1_160 ( .A(new_wire_519), .B(_265_), .C(_254_), .Y(AI_7_) );
INVX1 INVX1_104 ( .A(op_0_), .Y(_266_) );
INVX1 INVX1_105 ( .A(new_wire_494), .Y(_267_) );
NOR3X1 NOR3X1_14 ( .A(_816_), .B(_1130_), .C(new_wire_494), .Y(_268_) );
INVX2 INVX2_36 ( .A(new_wire_510), .Y(_269_) );
OAI21X1 OAI21X1_161 ( .A(new_wire_30), .B(new_wire_340), .C(new_wire_522), .Y(_270_) );
NOR2X1 NOR2X1_144 ( .A(_270_), .B(_121_), .Y(_271_) );
NAND2X1 NAND2X1_142 ( .A(new_wire_206), .B(_271_), .Y(_272_) );
NOR2X1 NOR2X1_145 ( .A(_268_), .B(_272_), .Y(_273_) );
OAI21X1 OAI21X1_162 ( .A(_266_), .B(_267_), .C(_273_), .Y(alu_op_0_) );
INVX1 INVX1_106 ( .A(op_1_), .Y(_274_) );
OAI21X1 OAI21X1_163 ( .A(_274_), .B(_267_), .C(_273_), .Y(alu_op_1_) );
INVX1 INVX1_107 ( .A(backwards), .Y(_275_) );
INVX1 INVX1_108 ( .A(_271_), .Y(_276_) );
AOI21X1 AOI21X1_60 ( .A(op_2_), .B(new_wire_494), .C(_276_), .Y(_277_) );
OAI21X1 OAI21X1_164 ( .A(_275_), .B(new_wire_208), .C(_277_), .Y(alu_op_2_) );
INVX1 INVX1_109 ( .A(op_3_), .Y(_278_) );
NOR2X1 NOR2X1_146 ( .A(_278_), .B(_267_), .Y(alu_op_3_) );
INVX1 INVX1_110 ( .A(store), .Y(_279_) );
OAI21X1 OAI21X1_165 ( .A(new_wire_33), .B(new_wire_432), .C(_271_), .Y(_280_) );
INVX1 INVX1_111 ( .A(new_wire_534), .Y(_281_) );
AND2X2 AND2X2_35 ( .A(_1199_), .B(_1190_), .Y(_282_) );
OAI21X1 OAI21X1_166 ( .A(_279_), .B(_282_), .C(_281_), .Y(_1441_) );
INVX2 INVX2_37 ( .A(new_wire_447), .Y(_283_) );
MUX2X1 MUX2X1_10 ( .A(C), .B(new_wire_331), .S(php), .Y(_284_) );
OAI22X1 OAI22X1_28 ( .A(_79_), .B(new_wire_270), .C(_284_), .D(new_wire_500), .Y(_285_) );
AOI21X1 AOI21X1_61 ( .A(new_wire_331), .B(new_wire_537), .C(_285_), .Y(_286_) );
INVX2 INVX2_38 ( .A(new_wire_498), .Y(_287_) );
AOI22X1 AOI22X1_26 ( .A(PC_8_), .B(new_wire_510), .C(PC_0_), .D(new_wire_539), .Y(_288_) );
AND2X2 AND2X2_36 ( .A(_286_), .B(_288_), .Y(_289_) );
OAI21X1 OAI21X1_167 ( .A(new_wire_534), .B(_163_), .C(_289_), .Y(_1440__0_) );
INVX1 INVX1_112 ( .A(php), .Y(_290_) );
OAI21X1 OAI21X1_168 ( .A(_290_), .B(new_wire_500), .C(new_wire_270), .Y(_291_) );
AOI22X1 AOI22X1_27 ( .A(PC_9_), .B(new_wire_510), .C(PC_1_), .D(new_wire_539), .Y(_292_) );
OAI21X1 OAI21X1_169 ( .A(php), .B(new_wire_500), .C(new_wire_447), .Y(_293_) );
INVX1 INVX1_113 ( .A(new_wire_541), .Y(_294_) );
OAI21X1 OAI21X1_170 ( .A(new_wire_347), .B(_294_), .C(_292_), .Y(_295_) );
AOI21X1 AOI21X1_62 ( .A(Z), .B(_291_), .C(_295_), .Y(_296_) );
OAI21X1 OAI21X1_171 ( .A(new_wire_534), .B(_186_), .C(_296_), .Y(_1440__1_) );
NAND2X1 NAND2X1_143 ( .A(new_wire_357), .B(new_wire_541), .Y(_297_) );
OAI22X1 OAI22X1_29 ( .A(new_wire_370), .B(new_wire_522), .C(new_wire_360), .D(new_wire_498), .Y(_298_) );
AOI21X1 AOI21X1_63 ( .A(I), .B(_291_), .C(_298_), .Y(_299_) );
AND2X2 AND2X2_37 ( .A(_299_), .B(_297_), .Y(_300_) );
OAI21X1 OAI21X1_172 ( .A(new_wire_534), .B(_199_), .C(_300_), .Y(_1440__2_) );
NOR2X1 NOR2X1_147 ( .A(_290_), .B(new_wire_501), .Y(_301_) );
OAI21X1 OAI21X1_173 ( .A(new_wire_304), .B(_301_), .C(new_wire_543), .Y(_302_) );
OAI22X1 OAI22X1_30 ( .A(new_wire_364), .B(new_wire_522), .C(new_wire_354), .D(new_wire_499), .Y(_303_) );
AOI21X1 AOI21X1_64 ( .A(new_wire_352), .B(new_wire_541), .C(_303_), .Y(_304_) );
AND2X2 AND2X2_38 ( .A(_304_), .B(_302_), .Y(_305_) );
OAI21X1 OAI21X1_174 ( .A(new_wire_535), .B(_212_), .C(_305_), .Y(_1440__3_) );
OAI22X1 OAI22X1_31 ( .A(new_wire_537), .B(new_wire_484), .C(new_wire_313), .D(_301_), .Y(_306_) );
OAI21X1 OAI21X1_175 ( .A(new_wire_271), .B(_829_), .C(_306_), .Y(_307_) );
OAI22X1 OAI22X1_32 ( .A(new_wire_376), .B(new_wire_522), .C(new_wire_318), .D(new_wire_499), .Y(_308_) );
NOR2X1 NOR2X1_148 ( .A(_308_), .B(_307_), .Y(_309_) );
OAI21X1 OAI21X1_176 ( .A(new_wire_535), .B(_225_), .C(_309_), .Y(_1440__4_) );
OAI22X1 OAI22X1_33 ( .A(new_wire_537), .B(new_wire_485), .C(new_wire_296), .D(_301_), .Y(_310_) );
OAI21X1 OAI21X1_177 ( .A(_787_), .B(new_wire_523), .C(new_wire_271), .Y(_311_) );
AOI21X1 AOI21X1_65 ( .A(PC_5_), .B(new_wire_539), .C(_311_), .Y(_312_) );
AND2X2 AND2X2_39 ( .A(_312_), .B(_310_), .Y(_313_) );
OAI21X1 OAI21X1_178 ( .A(new_wire_535), .B(_239_), .C(_313_), .Y(_1440__5_) );
INVX1 INVX1_114 ( .A(_291_), .Y(_314_) );
AOI22X1 AOI22X1_28 ( .A(PC_14_), .B(new_wire_511), .C(PC_6_), .D(new_wire_539), .Y(_315_) );
OAI21X1 OAI21X1_179 ( .A(_1306_), .B(_314_), .C(_315_), .Y(_316_) );
AOI21X1 AOI21X1_66 ( .A(new_wire_326), .B(new_wire_541), .C(_316_), .Y(_317_) );
OAI21X1 OAI21X1_180 ( .A(new_wire_535), .B(_252_), .C(_317_), .Y(_1440__6_) );
INVX1 INVX1_115 ( .A(N), .Y(_318_) );
AOI22X1 AOI22X1_29 ( .A(PC_15_), .B(new_wire_511), .C(PC_7_), .D(new_wire_540), .Y(_319_) );
OAI21X1 OAI21X1_181 ( .A(_318_), .B(_314_), .C(_319_), .Y(_320_) );
AOI21X1 AOI21X1_67 ( .A(new_wire_321), .B(new_wire_542), .C(_320_), .Y(_321_) );
OAI21X1 OAI21X1_182 ( .A(new_wire_536), .B(_265_), .C(_321_), .Y(_1440__7_) );
AND2X2 AND2X2_40 ( .A(new_wire_543), .B(adc_sbc), .Y(_14_) );
INVX1 INVX1_116 ( .A(adc_bcd), .Y(_322_) );
NOR2X1 NOR2X1_149 ( .A(_322_), .B(new_wire_452), .Y(ALU_BCD) );
INVX4 INVX4_6 ( .A(reset), .Y(_1175_) );
INVX1 INVX1_117 ( .A(res), .Y(_323_) );
OAI21X1 OAI21X1_183 ( .A(_323_), .B(_859__bF_buf0), .C(new_wire_545), .Y(_31_) );
INVX2 INVX2_39 ( .A(new_wire_547), .Y(_324_) );
NOR2X1 NOR2X1_150 ( .A(new_wire_549), .B(new_wire_119), .Y(_325_) );
OAI21X1 OAI21X1_184 ( .A(_828_), .B(_325_), .C(_169_), .Y(_326_) );
AOI21X1 AOI21X1_68 ( .A(new_wire_357), .B(_325_), .C(_326_), .Y(_327_) );
INVX1 INVX1_118 ( .A(new_wire_342), .Y(_328_) );
AOI21X1 AOI21X1_69 ( .A(new_wire_434), .B(new_wire_368), .C(_328_), .Y(_329_) );
INVX2 INVX2_40 ( .A(new_wire_434), .Y(_330_) );
INVX1 INVX1_119 ( .A(sei), .Y(_331_) );
AOI21X1 AOI21X1_70 ( .A(_828_), .B(_331_), .C(cli), .Y(_332_) );
OAI21X1 OAI21X1_185 ( .A(_332_), .B(_169_), .C(new_wire_551), .Y(_333_) );
OAI21X1 OAI21X1_186 ( .A(_333_), .B(_327_), .C(_329_), .Y(_6_) );
AND2X2 AND2X2_41 ( .A(new_wire_495), .B(shift_right), .Y(alu_shift_right) );
OAI21X1 OAI21X1_187 ( .A(_811_), .B(new_wire_132), .C(new_wire_342), .Y(_334_) );
OAI21X1 OAI21X1_188 ( .A(new_wire_132), .B(new_wire_439), .C(_136_), .Y(_335_) );
NOR2X1 NOR2X1_151 ( .A(_334_), .B(_335_), .Y(_336_) );
OAI21X1 OAI21X1_189 ( .A(new_wire_30), .B(new_wire_426), .C(_1201_), .Y(_337_) );
INVX1 INVX1_120 ( .A(load_reg), .Y(_338_) );
NOR2X1 NOR2X1_152 ( .A(new_wire_547), .B(_338_), .Y(_339_) );
AOI21X1 AOI21X1_71 ( .A(new_wire_197), .B(_339_), .C(_337_), .Y(_340_) );
AOI21X1 AOI21X1_72 ( .A(_336_), .B(_340_), .C(new_wire_190), .Y(_341_) );
NAND3X1 NAND3X1_131 ( .A(new_wire_127), .B(_341_), .C(new_wire_202), .Y(_342_) );
NOR2X1 NOR2X1_153 ( .A(new_wire_514), .B(_342_), .Y(_343_) );
OAI21X1 OAI21X1_190 ( .A(new_wire_132), .B(new_wire_439), .C(_904_), .Y(_344_) );
OAI21X1 OAI21X1_191 ( .A(new_wire_375), .B(new_wire_492), .C(_344_), .Y(_345_) );
MUX2X1 MUX2X1_11 ( .A(_345_), .B(_147_), .S(new_wire_557), .Y(_1442__0_) );
NOR2X1 NOR2X1_154 ( .A(adc_bcd), .B(HC), .Y(_346_) );
NAND2X1 NAND2X1_144 ( .A(adj_bcd), .B(_346_), .Y(_347_) );
NAND3X1 NAND3X1_132 ( .A(adc_bcd), .B(adj_bcd), .C(HC), .Y(_348_) );
NAND2X1 NAND2X1_145 ( .A(_348_), .B(_347_), .Y(_349_) );
INVX1 INVX1_121 ( .A(_349_), .Y(_350_) );
NAND2X1 NAND2X1_146 ( .A(new_wire_347), .B(_350_), .Y(_351_) );
NOR2X1 NOR2X1_155 ( .A(new_wire_347), .B(_350_), .Y(_352_) );
NOR2X1 NOR2X1_156 ( .A(new_wire_473), .B(_352_), .Y(_353_) );
AOI22X1 AOI22X1_30 ( .A(new_wire_372), .B(new_wire_474), .C(_351_), .D(_353_), .Y(_354_) );
MUX2X1 MUX2X1_12 ( .A(_354_), .B(_176_), .S(new_wire_557), .Y(_1442__1_) );
XNOR2X1 XNOR2X1_2 ( .A(_348_), .B(new_wire_357), .Y(_355_) );
INVX1 INVX1_122 ( .A(_355_), .Y(_356_) );
OAI21X1 OAI21X1_192 ( .A(new_wire_348), .B(_350_), .C(_356_), .Y(_357_) );
AOI21X1 AOI21X1_73 ( .A(_352_), .B(_355_), .C(new_wire_474), .Y(_358_) );
AOI22X1 AOI22X1_31 ( .A(new_wire_368), .B(new_wire_474), .C(_357_), .D(_358_), .Y(_359_) );
MUX2X1 MUX2X1_13 ( .A(_359_), .B(_189_), .S(new_wire_557), .Y(_1442__2_) );
INVX1 INVX1_123 ( .A(new_wire_358), .Y(_360_) );
NAND2X1 NAND2X1_147 ( .A(_355_), .B(_352_), .Y(_361_) );
OAI21X1 OAI21X1_193 ( .A(_360_), .B(_348_), .C(_361_), .Y(_362_) );
INVX2 INVX2_41 ( .A(new_wire_352), .Y(_363_) );
XNOR2X1 XNOR2X1_3 ( .A(_347_), .B(_363_), .Y(_364_) );
XNOR2X1 XNOR2X1_4 ( .A(_362_), .B(_364_), .Y(_365_) );
MUX2X1 MUX2X1_14 ( .A(_365_), .B(new_wire_362), .S(new_wire_492), .Y(_366_) );
MUX2X1 MUX2X1_15 ( .A(_366_), .B(_202_), .S(new_wire_557), .Y(_1442__3_) );
INVX1 INVX1_124 ( .A(new_wire_313), .Y(_367_) );
OAI21X1 OAI21X1_194 ( .A(new_wire_133), .B(new_wire_439), .C(_367_), .Y(_368_) );
OAI21X1 OAI21X1_195 ( .A(DIMUX_4_), .B(new_wire_492), .C(_368_), .Y(_369_) );
MUX2X1 MUX2X1_16 ( .A(_369_), .B(_215_), .S(new_wire_558), .Y(_1442__4_) );
INVX1 INVX1_125 ( .A(new_wire_335), .Y(_370_) );
NAND3X1 NAND3X1_133 ( .A(adj_bcd), .B(_370_), .C(_322_), .Y(_371_) );
NAND3X1 NAND3X1_134 ( .A(new_wire_336), .B(adc_bcd), .C(adj_bcd), .Y(_372_) );
NAND2X1 NAND2X1_148 ( .A(_372_), .B(_371_), .Y(_373_) );
INVX1 INVX1_126 ( .A(_373_), .Y(_374_) );
NAND2X1 NAND2X1_149 ( .A(new_wire_298), .B(_374_), .Y(_375_) );
NOR2X1 NOR2X1_157 ( .A(new_wire_298), .B(_374_), .Y(_376_) );
NOR2X1 NOR2X1_158 ( .A(new_wire_474), .B(_376_), .Y(_377_) );
AOI22X1 AOI22X1_32 ( .A(new_wire_293), .B(new_wire_475), .C(_375_), .D(_377_), .Y(_378_) );
MUX2X1 MUX2X1_17 ( .A(_378_), .B(_229_), .S(new_wire_558), .Y(_1442__5_) );
XNOR2X1 XNOR2X1_5 ( .A(_372_), .B(new_wire_326), .Y(_379_) );
INVX1 INVX1_127 ( .A(_379_), .Y(_380_) );
OAI21X1 OAI21X1_196 ( .A(new_wire_298), .B(_374_), .C(_380_), .Y(_381_) );
AOI21X1 AOI21X1_74 ( .A(_376_), .B(_379_), .C(new_wire_475), .Y(_382_) );
AOI22X1 AOI22X1_33 ( .A(new_wire_384), .B(new_wire_475), .C(_381_), .D(_382_), .Y(_383_) );
MUX2X1 MUX2X1_18 ( .A(_383_), .B(_242_), .S(new_wire_558), .Y(_1442__6_) );
INVX1 INVX1_128 ( .A(new_wire_326), .Y(_384_) );
NAND2X1 NAND2X1_150 ( .A(_379_), .B(_376_), .Y(_385_) );
OAI21X1 OAI21X1_197 ( .A(_384_), .B(_372_), .C(_385_), .Y(_386_) );
INVX2 INVX2_42 ( .A(new_wire_321), .Y(_387_) );
XNOR2X1 XNOR2X1_6 ( .A(_371_), .B(_387_), .Y(_388_) );
XNOR2X1 XNOR2X1_7 ( .A(_386_), .B(_388_), .Y(_389_) );
MUX2X1 MUX2X1_19 ( .A(_389_), .B(new_wire_388), .S(new_wire_493), .Y(_390_) );
MUX2X1 MUX2X1_20 ( .A(_390_), .B(_255_), .S(new_wire_558), .Y(_1442__7_) );
INVX1 INVX1_129 ( .A(NMI_1), .Y(_391_) );
NAND3X1 NAND3X1_135 ( .A(NMI), .B(new_wire_282), .C(_391_), .Y(_392_) );
OAI21X1 OAI21X1_198 ( .A(new_wire_282), .B(_328_), .C(_392_), .Y(_7_) );
NAND2X1 NAND2X1_151 ( .A(cond_code_0_), .B(new_wire_187), .Y(_393_) );
OAI21X1 OAI21X1_199 ( .A(new_wire_187), .B(_1361_), .C(_393_), .Y(_22__0_) );
NAND2X1 NAND2X1_152 ( .A(new_wire_483), .B(new_wire_177), .Y(_394_) );
OAI21X1 OAI21X1_200 ( .A(new_wire_177), .B(new_wire_453), .C(_394_), .Y(_22__1_) );
NAND2X1 NAND2X1_153 ( .A(cond_code_2_), .B(new_wire_177), .Y(_395_) );
OAI21X1 OAI21X1_201 ( .A(new_wire_178), .B(new_wire_408), .C(_395_), .Y(_22__2_) );
NAND2X1 NAND2X1_154 ( .A(new_wire_162), .B(new_wire_461), .Y(_396_) );
OAI22X1 OAI22X1_34 ( .A(new_wire_549), .B(new_wire_158), .C(new_wire_476), .D(_396_), .Y(_30_) );
INVX1 INVX1_130 ( .A(_1097_), .Y(_397_) );
NOR2X1 NOR2X1_159 ( .A(new_wire_80), .B(new_wire_467), .Y(_398_) );
INVX1 INVX1_131 ( .A(_398_), .Y(_399_) );
OAI22X1 OAI22X1_35 ( .A(_290_), .B(new_wire_158), .C(_399_), .D(_397_), .Y(_29_) );
OAI21X1 OAI21X1_202 ( .A(new_wire_187), .B(new_wire_120), .C(clc), .Y(_400_) );
OAI21X1 OAI21X1_203 ( .A(new_wire_106), .B(new_wire_413), .C(new_wire_423), .Y(_401_) );
NAND3X1 NAND3X1_136 ( .A(new_wire_408), .B(_398_), .C(new_wire_461), .Y(_402_) );
OAI21X1 OAI21X1_204 ( .A(_401_), .B(_402_), .C(_400_), .Y(_17_) );
OAI21X1 OAI21X1_205 ( .A(new_wire_191), .B(new_wire_114), .C(sec), .Y(_403_) );
NOR2X1 NOR2X1_160 ( .A(new_wire_442), .B(_1361_), .Y(_404_) );
INVX1 INVX1_132 ( .A(_404_), .Y(_405_) );
OAI21X1 OAI21X1_206 ( .A(_405_), .B(_402_), .C(_403_), .Y(_33_) );
OAI21X1 OAI21X1_207 ( .A(new_wire_188), .B(new_wire_120), .C(cld), .Y(_406_) );
OR2X2 OR2X2_18 ( .A(_401_), .B(new_wire_82), .Y(_407_) );
NOR2X1 NOR2X1_161 ( .A(new_wire_408), .B(new_wire_453), .Y(_408_) );
NAND2X1 NAND2X1_155 ( .A(_408_), .B(new_wire_462), .Y(_409_) );
OAI21X1 OAI21X1_208 ( .A(_407_), .B(_409_), .C(_406_), .Y(_18_) );
OAI21X1 OAI21X1_209 ( .A(new_wire_188), .B(new_wire_120), .C(sed), .Y(_410_) );
NAND2X1 NAND2X1_156 ( .A(new_wire_162), .B(_404_), .Y(_411_) );
OAI21X1 OAI21X1_210 ( .A(_411_), .B(_409_), .C(_410_), .Y(_34_) );
OAI21X1 OAI21X1_211 ( .A(new_wire_191), .B(new_wire_120), .C(cli), .Y(_412_) );
NOR2X1 NOR2X1_162 ( .A(new_wire_454), .B(new_wire_463), .Y(_413_) );
NAND2X1 NAND2X1_157 ( .A(_413_), .B(new_wire_462), .Y(_414_) );
OAI21X1 OAI21X1_212 ( .A(_407_), .B(_414_), .C(_412_), .Y(_19_) );
OAI22X1 OAI22X1_36 ( .A(_331_), .B(new_wire_162), .C(_411_), .D(_414_), .Y(_35_) );
NOR2X1 NOR2X1_163 ( .A(new_wire_408), .B(new_wire_467), .Y(_415_) );
NAND2X1 NAND2X1_158 ( .A(new_wire_559), .B(_404_), .Y(_416_) );
OAI21X1 OAI21X1_213 ( .A(new_wire_188), .B(new_wire_122), .C(clv), .Y(_417_) );
OAI21X1 OAI21X1_214 ( .A(_416_), .B(_396_), .C(_417_), .Y(_20_) );
OAI21X1 OAI21X1_215 ( .A(new_wire_101), .B(new_wire_402), .C(new_wire_399), .Y(_418_) );
INVX1 INVX1_133 ( .A(_418_), .Y(_419_) );
OAI21X1 OAI21X1_216 ( .A(new_wire_107), .B(_1082_), .C(_419_), .Y(_420_) );
OR2X2 OR2X2_19 ( .A(_420_), .B(new_wire_476), .Y(_421_) );
OAI21X1 OAI21X1_217 ( .A(new_wire_191), .B(new_wire_114), .C(bit_ins), .Y(_422_) );
OAI21X1 OAI21X1_218 ( .A(new_wire_78), .B(_421_), .C(_422_), .Y(_16_) );
NAND2X1 NAND2X1_159 ( .A(new_wire_409), .B(new_wire_488), .Y(_423_) );
INVX1 INVX1_134 ( .A(_408_), .Y(_424_) );
INVX1 INVX1_135 ( .A(new_wire_446), .Y(_425_) );
NOR2X1 NOR2X1_164 ( .A(new_wire_430), .B(new_wire_416), .Y(_426_) );
AOI21X1 AOI21X1_75 ( .A(new_wire_488), .B(_426_), .C(_425_), .Y(_427_) );
NAND3X1 NAND3X1_137 ( .A(new_wire_464), .B(_1095_), .C(new_wire_462), .Y(_428_) );
OAI22X1 OAI22X1_37 ( .A(_424_), .B(_427_), .C(new_wire_468), .D(_428_), .Y(_429_) );
NOR2X1 NOR2X1_165 ( .A(new_wire_460), .B(_424_), .Y(_430_) );
NOR2X1 NOR2X1_166 ( .A(new_wire_423), .B(_424_), .Y(_431_) );
AOI22X1 AOI22X1_34 ( .A(_430_), .B(_1136_), .C(new_wire_470), .D(_431_), .Y(_432_) );
NAND3X1 NAND3X1_138 ( .A(_1187_), .B(_1227_), .C(_1359_), .Y(_433_) );
NAND2X1 NAND2X1_160 ( .A(_433_), .B(_432_), .Y(_434_) );
NOR2X1 NOR2X1_167 ( .A(_429_), .B(_434_), .Y(_435_) );
NAND3X1 NAND3X1_139 ( .A(new_wire_409), .B(_1299_), .C(_425_), .Y(_436_) );
INVX1 INVX1_136 ( .A(_436_), .Y(_437_) );
NAND2X1 NAND2X1_161 ( .A(_413_), .B(new_wire_488), .Y(_438_) );
OAI21X1 OAI21X1_219 ( .A(new_wire_476), .B(_420_), .C(_438_), .Y(_439_) );
NOR2X1 NOR2X1_168 ( .A(_437_), .B(_439_), .Y(_440_) );
NAND2X1 NAND2X1_162 ( .A(_440_), .B(_435_), .Y(_441_) );
INVX1 INVX1_137 ( .A(_441_), .Y(_442_) );
OAI21X1 OAI21X1_220 ( .A(new_wire_468), .B(_423_), .C(_442_), .Y(_443_) );
INVX1 INVX1_138 ( .A(_435_), .Y(_444_) );
NOR2X1 NOR2X1_169 ( .A(new_wire_477), .B(_420_), .Y(_445_) );
OAI21X1 OAI21X1_221 ( .A(new_wire_464), .B(new_wire_486), .C(new_wire_160), .Y(_446_) );
NOR2X1 NOR2X1_170 ( .A(_446_), .B(_445_), .Y(_447_) );
OAI21X1 OAI21X1_222 ( .A(_1361_), .B(_436_), .C(_447_), .Y(_448_) );
NOR2X1 NOR2X1_171 ( .A(_448_), .B(_444_), .Y(_449_) );
AOI22X1 AOI22X1_35 ( .A(_266_), .B(new_wire_78), .C(_449_), .D(_443_), .Y(_28__0_) );
NOR2X1 NOR2X1_172 ( .A(_1276_), .B(new_wire_446), .Y(_450_) );
AOI21X1 AOI21X1_76 ( .A(_450_), .B(new_wire_409), .C(_446_), .Y(_451_) );
AND2X2 AND2X2_42 ( .A(_435_), .B(_451_), .Y(_452_) );
AOI22X1 AOI22X1_36 ( .A(_274_), .B(new_wire_78), .C(_441_), .D(_452_), .Y(_28__1_) );
OAI21X1 OAI21X1_223 ( .A(new_wire_191), .B(new_wire_114), .C(op_2_), .Y(_453_) );
OAI21X1 OAI21X1_224 ( .A(new_wire_78), .B(_442_), .C(_453_), .Y(_28__2_) );
AOI22X1 AOI22X1_37 ( .A(_278_), .B(new_wire_79), .C(_436_), .D(_447_), .Y(_28__3_) );
NAND3X1 NAND3X1_140 ( .A(_1083_), .B(new_wire_416), .C(_419_), .Y(_454_) );
NOR2X1 NOR2X1_173 ( .A(new_wire_464), .B(_454_), .Y(_455_) );
AOI21X1 AOI21X1_77 ( .A(_1362_), .B(_1359_), .C(_455_), .Y(_456_) );
OAI21X1 OAI21X1_225 ( .A(new_wire_192), .B(new_wire_122), .C(rotate), .Y(_457_) );
OAI21X1 OAI21X1_226 ( .A(new_wire_82), .B(_456_), .C(_457_), .Y(_32_) );
OAI21X1 OAI21X1_227 ( .A(new_wire_192), .B(new_wire_114), .C(shift_right), .Y(_458_) );
OAI21X1 OAI21X1_228 ( .A(new_wire_79), .B(_438_), .C(_458_), .Y(_37_) );
AOI21X1 AOI21X1_78 ( .A(_450_), .B(new_wire_464), .C(new_wire_82), .Y(_459_) );
AOI22X1 AOI22X1_38 ( .A(new_wire_496), .B(new_wire_82), .C(_459_), .D(_432_), .Y(_21_) );
OAI21X1 OAI21X1_229 ( .A(new_wire_399), .B(_1181_), .C(new_wire_160), .Y(_460_) );
OAI22X1 OAI22X1_38 ( .A(_87_), .B(new_wire_162), .C(_460_), .D(_423_), .Y(_36_) );
OAI21X1 OAI21X1_230 ( .A(new_wire_197), .B(_1123_), .C(new_wire_26), .Y(_461_) );
INVX1 INVX1_139 ( .A(_461_), .Y(_462_) );
NAND2X1 NAND2X1_163 ( .A(new_wire_543), .B(new_wire_409), .Y(_463_) );
NOR2X1 NOR2X1_174 ( .A(_1299_), .B(new_wire_446), .Y(_464_) );
NAND2X1 NAND2X1_164 ( .A(_462_), .B(_464_), .Y(_465_) );
OAI22X1 OAI22X1_39 ( .A(_322_), .B(_462_), .C(_463_), .D(_465_), .Y(_12_) );
INVX2 INVX2_43 ( .A(adc_sbc), .Y(_466_) );
OAI21X1 OAI21X1_231 ( .A(_466_), .B(_462_), .C(_465_), .Y(_13_) );
OAI21X1 OAI21X1_232 ( .A(new_wire_424), .B(new_wire_405), .C(_454_), .Y(_467_) );
NAND2X1 NAND2X1_165 ( .A(_408_), .B(_467_), .Y(_468_) );
OAI21X1 OAI21X1_233 ( .A(new_wire_192), .B(new_wire_123), .C(inc), .Y(_469_) );
OAI21X1 OAI21X1_234 ( .A(new_wire_83), .B(_468_), .C(_469_), .Y(_24_) );
AND2X2 AND2X2_43 ( .A(new_wire_111), .B(_341_), .Y(_470_) );
NAND2X1 NAND2X1_166 ( .A(new_wire_517), .B(_470_), .Y(_471_) );
NAND2X1 NAND2X1_167 ( .A(AXYS_0__0_), .B(new_wire_561), .Y(_472_) );
OAI21X1 OAI21X1_235 ( .A(_345_), .B(new_wire_561), .C(_472_), .Y(_1443__0_) );
NAND2X1 NAND2X1_168 ( .A(AXYS_0__1_), .B(new_wire_561), .Y(_473_) );
OAI21X1 OAI21X1_236 ( .A(_354_), .B(new_wire_561), .C(_473_), .Y(_1443__1_) );
NAND2X1 NAND2X1_169 ( .A(AXYS_0__2_), .B(new_wire_562), .Y(_474_) );
OAI21X1 OAI21X1_237 ( .A(_359_), .B(new_wire_562), .C(_474_), .Y(_1443__2_) );
NAND2X1 NAND2X1_170 ( .A(AXYS_0__3_), .B(new_wire_562), .Y(_475_) );
OAI21X1 OAI21X1_238 ( .A(_366_), .B(new_wire_562), .C(_475_), .Y(_1443__3_) );
NAND2X1 NAND2X1_171 ( .A(AXYS_0__4_), .B(new_wire_563), .Y(_476_) );
OAI21X1 OAI21X1_239 ( .A(_369_), .B(new_wire_563), .C(_476_), .Y(_1443__4_) );
NAND2X1 NAND2X1_172 ( .A(AXYS_0__5_), .B(new_wire_563), .Y(_477_) );
OAI21X1 OAI21X1_240 ( .A(_378_), .B(new_wire_563), .C(_477_), .Y(_1443__5_) );
NAND2X1 NAND2X1_173 ( .A(AXYS_0__6_), .B(new_wire_564), .Y(_478_) );
OAI21X1 OAI21X1_241 ( .A(_383_), .B(new_wire_564), .C(_478_), .Y(_1443__6_) );
NAND2X1 NAND2X1_174 ( .A(AXYS_0__7_), .B(new_wire_564), .Y(_479_) );
OAI21X1 OAI21X1_242 ( .A(_390_), .B(new_wire_564), .C(_479_), .Y(_1443__7_) );
NAND2X1 NAND2X1_175 ( .A(new_wire_416), .B(new_wire_559), .Y(_480_) );
OAI21X1 OAI21X1_243 ( .A(new_wire_192), .B(new_wire_115), .C(load_only), .Y(_481_) );
OAI21X1 OAI21X1_244 ( .A(new_wire_83), .B(_480_), .C(_481_), .Y(_26_) );
INVX1 INVX1_140 ( .A(new_wire_559), .Y(_482_) );
NAND3X1 NAND3X1_141 ( .A(_1141_), .B(new_wire_489), .C(_482_), .Y(_483_) );
OAI21X1 OAI21X1_245 ( .A(_1212_), .B(new_wire_157), .C(_483_), .Y(_40_) );
NOR2X1 NOR2X1_175 ( .A(new_wire_410), .B(new_wire_417), .Y(_484_) );
OAI21X1 OAI21X1_246 ( .A(_419_), .B(_425_), .C(_484_), .Y(_485_) );
OAI22X1 OAI22X1_40 ( .A(_279_), .B(new_wire_158), .C(_399_), .D(_485_), .Y(_39_) );
NOR2X1 NOR2X1_176 ( .A(new_wire_487), .B(_482_), .Y(_486_) );
NAND3X1 NAND3X1_142 ( .A(new_wire_400), .B(_1331_), .C(_486_), .Y(_487_) );
MUX2X1 MUX2X1_21 ( .A(_1184_), .B(index_y), .S(new_wire_155), .Y(_488_) );
NAND3X1 NAND3X1_143 ( .A(_1322_), .B(_488_), .C(_487_), .Y(_25_) );
INVX1 INVX1_141 ( .A(src_reg_0_), .Y(_489_) );
NAND3X1 NAND3X1_144 ( .A(new_wire_559), .B(_426_), .C(new_wire_403), .Y(_490_) );
NOR2X1 NOR2X1_177 ( .A(_401_), .B(_482_), .Y(_491_) );
INVX1 INVX1_142 ( .A(_491_), .Y(_492_) );
OAI21X1 OAI21X1_247 ( .A(new_wire_406), .B(_492_), .C(_490_), .Y(_493_) );
OAI21X1 OAI21X1_248 ( .A(new_wire_107), .B(new_wire_414), .C(new_wire_442), .Y(_494_) );
INVX1 INVX1_143 ( .A(_430_), .Y(_495_) );
OAI21X1 OAI21X1_249 ( .A(_494_), .B(_495_), .C(_428_), .Y(_496_) );
NOR2X1 NOR2X1_178 ( .A(_496_), .B(_493_), .Y(_497_) );
OAI21X1 OAI21X1_250 ( .A(new_wire_490), .B(_416_), .C(_497_), .Y(_498_) );
NAND2X1 NAND2X1_176 ( .A(new_wire_158), .B(_498_), .Y(_499_) );
OAI21X1 OAI21X1_251 ( .A(_489_), .B(new_wire_159), .C(_499_), .Y(_38__0_) );
NAND2X1 NAND2X1_177 ( .A(_408_), .B(_1095_), .Y(_500_) );
OAI21X1 OAI21X1_252 ( .A(_500_), .B(new_wire_490), .C(new_wire_161), .Y(_501_) );
NOR2X1 NOR2X1_179 ( .A(new_wire_417), .B(_1077_), .Y(_502_) );
OAI21X1 OAI21X1_253 ( .A(_426_), .B(_502_), .C(_486_), .Y(_503_) );
OAI21X1 OAI21X1_254 ( .A(_1268_), .B(_495_), .C(_503_), .Y(_504_) );
NOR2X1 NOR2X1_180 ( .A(_501_), .B(_504_), .Y(_505_) );
AOI22X1 AOI22X1_39 ( .A(_128_), .B(new_wire_81), .C(_505_), .D(_497_), .Y(_38__1_) );
INVX1 INVX1_144 ( .A(dst_reg_0_), .Y(_506_) );
OAI21X1 OAI21X1_255 ( .A(new_wire_442), .B(new_wire_400), .C(new_wire_404), .Y(_507_) );
OAI21X1 OAI21X1_256 ( .A(_480_), .B(_507_), .C(_428_), .Y(_508_) );
OAI21X1 OAI21X1_257 ( .A(new_wire_490), .B(_492_), .C(_397_), .Y(_509_) );
OAI21X1 OAI21X1_258 ( .A(_508_), .B(_509_), .C(new_wire_163), .Y(_510_) );
OAI21X1 OAI21X1_259 ( .A(_506_), .B(new_wire_159), .C(_510_), .Y(_23__0_) );
AOI21X1 AOI21X1_79 ( .A(new_wire_417), .B(_486_), .C(_501_), .Y(_511_) );
OAI21X1 OAI21X1_260 ( .A(_1268_), .B(_409_), .C(_511_), .Y(_512_) );
NOR2X1 NOR2X1_181 ( .A(_508_), .B(_512_), .Y(_513_) );
AOI21X1 AOI21X1_80 ( .A(_141_), .B(new_wire_81), .C(_513_), .Y(_23__1_) );
OAI21X1 OAI21X1_261 ( .A(new_wire_491), .B(_416_), .C(_433_), .Y(_514_) );
NOR2X1 NOR2X1_182 ( .A(_418_), .B(_416_), .Y(_515_) );
NOR2X1 NOR2X1_183 ( .A(new_wire_400), .B(_1085_), .Y(_516_) );
NAND3X1 NAND3X1_145 ( .A(_516_), .B(new_wire_560), .C(_502_), .Y(_517_) );
OAI21X1 OAI21X1_262 ( .A(new_wire_466), .B(new_wire_491), .C(_517_), .Y(_518_) );
NOR2X1 NOR2X1_184 ( .A(_515_), .B(_518_), .Y(_519_) );
OAI21X1 OAI21X1_263 ( .A(_1188_), .B(_1292_), .C(_519_), .Y(_520_) );
OAI22X1 OAI22X1_41 ( .A(new_wire_446), .B(_484_), .C(new_wire_424), .D(new_wire_406), .Y(_521_) );
OR2X2 OR2X2_20 ( .A(_520_), .B(_521_), .Y(_522_) );
OAI21X1 OAI21X1_264 ( .A(_514_), .B(_522_), .C(new_wire_161), .Y(_523_) );
OAI21X1 OAI21X1_265 ( .A(_338_), .B(new_wire_157), .C(_523_), .Y(_27_) );
OAI21X1 OAI21X1_266 ( .A(new_wire_392), .B(new_wire_458), .C(new_wire_26), .Y(_524_) );
OR2X2 OR2X2_21 ( .A(new_wire_565), .B(reset), .Y(_525_) );
OAI21X1 OAI21X1_267 ( .A(reset), .B(new_wire_565), .C(IRHOLD_0_), .Y(_526_) );
OAI21X1 OAI21X1_268 ( .A(_104_), .B(new_wire_567), .C(_526_), .Y(_4__0_) );
OAI21X1 OAI21X1_269 ( .A(reset), .B(new_wire_565), .C(IRHOLD_1_), .Y(_527_) );
OAI21X1 OAI21X1_270 ( .A(_118_), .B(new_wire_567), .C(_527_), .Y(_4__1_) );
OAI21X1 OAI21X1_271 ( .A(reset), .B(new_wire_565), .C(IRHOLD_2_), .Y(_528_) );
OAI21X1 OAI21X1_272 ( .A(new_wire_367), .B(new_wire_567), .C(_528_), .Y(_4__2_) );
OAI21X1 OAI21X1_273 ( .A(reset), .B(new_wire_566), .C(IRHOLD_3_), .Y(_529_) );
OAI21X1 OAI21X1_274 ( .A(_1179_), .B(new_wire_567), .C(_529_), .Y(_4__3_) );
INVX1 INVX1_145 ( .A(IRHOLD_4_), .Y(_530_) );
MUX2X1 MUX2X1_22 ( .A(_530_), .B(new_wire_379), .S(new_wire_568), .Y(_4__4_) );
INVX1 INVX1_146 ( .A(IRHOLD_5_), .Y(_531_) );
MUX2X1 MUX2X1_23 ( .A(_531_), .B(_119_), .S(new_wire_568), .Y(_4__5_) );
INVX1 INVX1_147 ( .A(IRHOLD_6_), .Y(_532_) );
MUX2X1 MUX2X1_24 ( .A(_532_), .B(new_wire_383), .S(new_wire_568), .Y(_4__6_) );
INVX1 INVX1_148 ( .A(IRHOLD_7_), .Y(_533_) );
MUX2X1 MUX2X1_25 ( .A(_533_), .B(new_wire_387), .S(new_wire_568), .Y(_4__7_) );
OAI21X1 OAI21X1_275 ( .A(new_wire_188), .B(new_wire_121), .C(new_wire_396), .Y(_534_) );
OAI21X1 OAI21X1_276 ( .A(reset), .B(_534_), .C(new_wire_569), .Y(_5_) );
AOI21X1 AOI21X1_81 ( .A(_1306_), .B(_466_), .C(new_wire_547), .Y(_535_) );
OAI21X1 OAI21X1_277 ( .A(_466_), .B(AV), .C(_535_), .Y(_536_) );
NOR2X1 NOR2X1_185 ( .A(clv), .B(_536_), .Y(_537_) );
AOI21X1 AOI21X1_82 ( .A(new_wire_326), .B(new_wire_547), .C(_537_), .Y(_538_) );
INVX1 INVX1_149 ( .A(bit_ins), .Y(_539_) );
NOR2X1 NOR2X1_186 ( .A(_539_), .B(new_wire_452), .Y(_540_) );
NAND2X1 NAND2X1_178 ( .A(new_wire_384), .B(_540_), .Y(_541_) );
OAI21X1 OAI21X1_278 ( .A(_1306_), .B(_540_), .C(_541_), .Y(_542_) );
NOR2X1 NOR2X1_187 ( .A(new_wire_198), .B(new_wire_434), .Y(_543_) );
AOI22X1 AOI22X1_40 ( .A(new_wire_384), .B(new_wire_435), .C(new_wire_570), .D(_542_), .Y(_544_) );
OAI21X1 OAI21X1_279 ( .A(new_wire_116), .B(_538_), .C(_544_), .Y(_10_) );
NAND2X1 NAND2X1_179 ( .A(new_wire_363), .B(new_wire_435), .Y(_545_) );
NOR2X1 NOR2X1_188 ( .A(new_wire_548), .B(cld), .Y(_546_) );
OAI21X1 OAI21X1_280 ( .A(new_wire_543), .B(sed), .C(_546_), .Y(_547_) );
OAI21X1 OAI21X1_281 ( .A(_363_), .B(new_wire_549), .C(_547_), .Y(_548_) );
MUX2X1 MUX2X1_26 ( .A(new_wire_544), .B(_548_), .S(new_wire_116), .Y(_549_) );
OAI21X1 OAI21X1_282 ( .A(new_wire_435), .B(_549_), .C(_545_), .Y(_3_) );
NAND2X1 NAND2X1_180 ( .A(new_wire_514), .B(_470_), .Y(_550_) );
NAND2X1 NAND2X1_181 ( .A(AXYS_2__0_), .B(new_wire_572), .Y(_551_) );
OAI21X1 OAI21X1_283 ( .A(_345_), .B(new_wire_572), .C(_551_), .Y(_1444__0_) );
NAND2X1 NAND2X1_182 ( .A(AXYS_2__1_), .B(new_wire_572), .Y(_552_) );
OAI21X1 OAI21X1_284 ( .A(_354_), .B(new_wire_572), .C(_552_), .Y(_1444__1_) );
NAND2X1 NAND2X1_183 ( .A(AXYS_2__2_), .B(new_wire_573), .Y(_553_) );
OAI21X1 OAI21X1_285 ( .A(_359_), .B(new_wire_573), .C(_553_), .Y(_1444__2_) );
NAND2X1 NAND2X1_184 ( .A(AXYS_2__3_), .B(new_wire_573), .Y(_554_) );
OAI21X1 OAI21X1_286 ( .A(_366_), .B(new_wire_573), .C(_554_), .Y(_1444__3_) );
NAND2X1 NAND2X1_185 ( .A(AXYS_2__4_), .B(new_wire_574), .Y(_555_) );
OAI21X1 OAI21X1_287 ( .A(_369_), .B(new_wire_574), .C(_555_), .Y(_1444__4_) );
NAND2X1 NAND2X1_186 ( .A(AXYS_2__5_), .B(new_wire_574), .Y(_556_) );
OAI21X1 OAI21X1_288 ( .A(_378_), .B(new_wire_574), .C(_556_), .Y(_1444__5_) );
NAND2X1 NAND2X1_187 ( .A(AXYS_2__6_), .B(new_wire_575), .Y(_557_) );
OAI21X1 OAI21X1_289 ( .A(_383_), .B(new_wire_575), .C(_557_), .Y(_1444__6_) );
NAND2X1 NAND2X1_188 ( .A(AXYS_2__7_), .B(new_wire_575), .Y(_558_) );
OAI21X1 OAI21X1_290 ( .A(_390_), .B(new_wire_575), .C(_558_), .Y(_1444__7_) );
INVX1 INVX1_150 ( .A(AN), .Y(_559_) );
OAI21X1 OAI21X1_291 ( .A(new_wire_514), .B(_155__bF_buf0), .C(load_reg), .Y(_560_) );
AOI21X1 AOI21X1_83 ( .A(_560_), .B(new_wire_496), .C(_559_), .Y(_561_) );
NAND2X1 NAND2X1_189 ( .A(new_wire_496), .B(_560_), .Y(_562_) );
OAI21X1 OAI21X1_292 ( .A(_318_), .B(_562_), .C(new_wire_549), .Y(_563_) );
AOI21X1 AOI21X1_84 ( .A(_387_), .B(new_wire_548), .C(new_wire_116), .Y(_564_) );
OAI21X1 OAI21X1_293 ( .A(_561_), .B(_563_), .C(_564_), .Y(_565_) );
OAI21X1 OAI21X1_294 ( .A(_539_), .B(new_wire_452), .C(new_wire_551), .Y(_566_) );
NAND2X1 NAND2X1_190 ( .A(N), .B(new_wire_570), .Y(_567_) );
OAI21X1 OAI21X1_295 ( .A(_540_), .B(_567_), .C(new_wire_447), .Y(_568_) );
AOI21X1 AOI21X1_85 ( .A(new_wire_388), .B(_566_), .C(_568_), .Y(_569_) );
AOI22X1 AOI22X1_41 ( .A(_559_), .B(new_wire_537), .C(_569_), .D(_565_), .Y(_8_) );
INVX1 INVX1_151 ( .A(AZ), .Y(_570_) );
NAND3X1 NAND3X1_146 ( .A(new_wire_497), .B(_539_), .C(_560_), .Y(_571_) );
AND2X2 AND2X2_44 ( .A(_571_), .B(AZ), .Y(_572_) );
OAI21X1 OAI21X1_296 ( .A(_1303_), .B(_571_), .C(new_wire_550), .Y(_573_) );
AOI21X1 AOI21X1_86 ( .A(new_wire_348), .B(new_wire_548), .C(new_wire_116), .Y(_574_) );
OAI21X1 OAI21X1_297 ( .A(_572_), .B(_573_), .C(_574_), .Y(_575_) );
OAI21X1 OAI21X1_298 ( .A(_118_), .B(new_wire_551), .C(new_wire_448), .Y(_576_) );
AOI21X1 AOI21X1_87 ( .A(new_wire_570), .B(Z), .C(_576_), .Y(_577_) );
AOI22X1 AOI22X1_42 ( .A(_570_), .B(new_wire_538), .C(_577_), .D(_575_), .Y(_11_) );
NOR2X1 NOR2X1_189 ( .A(_87_), .B(new_wire_448), .Y(_578_) );
NAND3X1 NAND3X1_147 ( .A(new_wire_497), .B(_87_), .C(_466_), .Y(_579_) );
NOR2X1 NOR2X1_190 ( .A(new_wire_548), .B(clc), .Y(_580_) );
OAI21X1 OAI21X1_299 ( .A(C), .B(sec), .C(_580_), .Y(_581_) );
OAI21X1 OAI21X1_300 ( .A(_904_), .B(new_wire_550), .C(_581_), .Y(_582_) );
NOR2X1 NOR2X1_191 ( .A(write_back), .B(new_wire_117), .Y(_583_) );
OAI21X1 OAI21X1_301 ( .A(_579_), .B(_582_), .C(_583_), .Y(_584_) );
AOI21X1 AOI21X1_88 ( .A(_370_), .B(_579_), .C(_584_), .Y(_585_) );
OAI21X1 OAI21X1_302 ( .A(_79_), .B(_583_), .C(new_wire_551), .Y(_586_) );
OAI22X1 OAI22X1_42 ( .A(new_wire_375), .B(new_wire_552), .C(_586_), .D(_585_), .Y(_587_) );
NAND2X1 NAND2X1_191 ( .A(new_wire_336), .B(_578_), .Y(_588_) );
OAI21X1 OAI21X1_303 ( .A(_578_), .B(_587_), .C(_588_), .Y(_2_) );
NOR2X1 NOR2X1_192 ( .A(new_wire_517), .B(_342_), .Y(_589_) );
MUX2X1 MUX2X1_27 ( .A(_345_), .B(_158_), .S(new_wire_576), .Y(_1445__0_) );
MUX2X1 MUX2X1_28 ( .A(_354_), .B(_181_), .S(new_wire_576), .Y(_1445__1_) );
MUX2X1 MUX2X1_29 ( .A(_359_), .B(_194_), .S(new_wire_576), .Y(_1445__2_) );
MUX2X1 MUX2X1_30 ( .A(_366_), .B(_207_), .S(new_wire_576), .Y(_1445__3_) );
MUX2X1 MUX2X1_31 ( .A(_369_), .B(_220_), .S(new_wire_577), .Y(_1445__4_) );
MUX2X1 MUX2X1_32 ( .A(_378_), .B(_234_), .S(new_wire_577), .Y(_1445__5_) );
MUX2X1 MUX2X1_33 ( .A(_383_), .B(_247_), .S(new_wire_577), .Y(_1445__6_) );
MUX2X1 MUX2X1_34 ( .A(_390_), .B(_260_), .S(new_wire_577), .Y(_1445__7_) );
NAND2X1 NAND2X1_192 ( .A(new_wire_27), .B(DI[7]), .Y(_590_) );
OAI21X1 OAI21X1_304 ( .A(new_wire_27), .B(_275_), .C(_590_), .Y(_15_) );
NOR2X1 NOR2X1_193 ( .A(_95_), .B(_270_), .Y(_591_) );
AOI21X1 AOI21X1_89 ( .A(_157_), .B(_162_), .C(new_wire_578), .Y(_592_) );
NOR2X1 NOR2X1_194 ( .A(_337_), .B(_94_), .Y(_593_) );
NAND3X1 NAND3X1_148 ( .A(new_wire_552), .B(_136_), .C(_593_), .Y(_594_) );
NOR2X1 NOR2X1_195 ( .A(_121_), .B(_594_), .Y(_595_) );
OAI21X1 OAI21X1_305 ( .A(new_wire_225), .B(new_wire_391), .C(_1211_), .Y(_596_) );
OR2X2 OR2X2_22 ( .A(_596_), .B(_91_), .Y(_597_) );
NOR2X1 NOR2X1_196 ( .A(new_wire_250), .B(_911_), .Y(_598_) );
OAI21X1 OAI21X1_306 ( .A(new_wire_133), .B(new_wire_391), .C(_598_), .Y(_599_) );
NOR2X1 NOR2X1_197 ( .A(_597_), .B(_599_), .Y(_600_) );
OAI21X1 OAI21X1_307 ( .A(new_wire_226), .B(new_wire_428), .C(_1109_), .Y(_601_) );
OAI21X1 OAI21X1_308 ( .A(new_wire_139), .B(new_wire_456), .C(_1115_), .Y(_602_) );
NOR2X1 NOR2X1_198 ( .A(_602_), .B(_601_), .Y(_603_) );
NAND3X1 NAND3X1_149 ( .A(_603_), .B(new_wire_581), .C(_595_), .Y(_604_) );
OAI21X1 OAI21X1_309 ( .A(new_wire_31), .B(new_wire_433), .C(_80_), .Y(_605_) );
OR2X2 OR2X2_23 ( .A(new_wire_586), .B(new_wire_90), .Y(_606_) );
NAND2X1 NAND2X1_193 ( .A(new_wire_248), .B(new_wire_343), .Y(_607_) );
NAND3X1 NAND3X1_150 ( .A(new_wire_301), .B(_607_), .C(_1197_), .Y(_608_) );
OAI21X1 OAI21X1_310 ( .A(new_wire_31), .B(new_wire_428), .C(_1320_), .Y(_609_) );
NOR2X1 NOR2X1_199 ( .A(_608_), .B(new_wire_588), .Y(_610_) );
NAND2X1 NAND2X1_194 ( .A(_610_), .B(new_wire_578), .Y(_611_) );
OR2X2 OR2X2_24 ( .A(_611_), .B(_606_), .Y(_612_) );
OR2X2 OR2X2_25 ( .A(_612_), .B(new_wire_583), .Y(_613_) );
INVX1 INVX1_152 ( .A(ABL_0_), .Y(_614_) );
AOI22X1 AOI22X1_43 ( .A(new_wire_331), .B(new_wire_92), .C(new_wire_375), .D(new_wire_588), .Y(_615_) );
NOR2X1 NOR2X1_200 ( .A(_608_), .B(new_wire_586), .Y(_616_) );
OAI21X1 OAI21X1_311 ( .A(_614_), .B(new_wire_595), .C(_615_), .Y(_617_) );
AOI21X1 AOI21X1_90 ( .A(new_wire_583), .B(new_wire_331), .C(_617_), .Y(_618_) );
OAI21X1 OAI21X1_312 ( .A(new_wire_333), .B(new_wire_591), .C(_618_), .Y(_619_) );
OR2X2 OR2X2_26 ( .A(_619_), .B(_592_), .Y(_1439__0_) );
OAI21X1 OAI21X1_313 ( .A(new_wire_344), .B(new_wire_450), .C(new_wire_248), .Y(_620_) );
INVX1 INVX1_153 ( .A(_135_), .Y(_621_) );
NAND2X1 NAND2X1_195 ( .A(_621_), .B(new_wire_570), .Y(_622_) );
AOI21X1 AOI21X1_91 ( .A(new_wire_248), .B(new_wire_288), .C(_1312_), .Y(_623_) );
NAND3X1 NAND3X1_151 ( .A(_166_), .B(_623_), .C(_598_), .Y(_624_) );
NOR2X1 NOR2X1_201 ( .A(_622_), .B(_624_), .Y(_625_) );
OR2X2 OR2X2_27 ( .A(_922_), .B(new_wire_317), .Y(_626_) );
NAND2X1 NAND2X1_196 ( .A(_107_), .B(_164_), .Y(_627_) );
OR2X2 OR2X2_28 ( .A(_626_), .B(_627_), .Y(_628_) );
NOR2X1 NOR2X1_202 ( .A(_122_), .B(_628_), .Y(_629_) );
NAND3X1 NAND3X1_152 ( .A(_620_), .B(_625_), .C(_629_), .Y(_630_) );
NOR2X1 NOR2X1_203 ( .A(new_wire_260), .B(_96_), .Y(_631_) );
NAND3X1 NAND3X1_153 ( .A(_136_), .B(_620_), .C(new_wire_501), .Y(_632_) );
NOR2X1 NOR2X1_204 ( .A(_632_), .B(_108_), .Y(_633_) );
NOR2X1 NOR2X1_205 ( .A(_328_), .B(new_wire_393), .Y(_634_) );
OAI21X1 OAI21X1_314 ( .A(_621_), .B(_634_), .C(new_wire_571), .Y(_635_) );
NOR2X1 NOR2X1_206 ( .A(_1336_), .B(_1099_), .Y(_636_) );
NOR2X1 NOR2X1_207 ( .A(_1416_), .B(new_wire_475), .Y(_637_) );
NAND3X1 NAND3X1_154 ( .A(_110_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_208 ( .A(_635_), .B(_638_), .Y(_639_) );
NAND3X1 NAND3X1_155 ( .A(_631_), .B(_633_), .C(_639_), .Y(_640_) );
NOR2X1 NOR2X1_209 ( .A(_596_), .B(_601_), .Y(_641_) );
NOR2X1 NOR2X1_210 ( .A(_337_), .B(new_wire_588), .Y(_642_) );
AND2X2 AND2X2_45 ( .A(_642_), .B(_641_), .Y(_643_) );
NAND3X1 NAND3X1_156 ( .A(_1197_), .B(_1115_), .C(_1150_), .Y(_644_) );
NAND3X1 NAND3X1_157 ( .A(_925_), .B(_1114_), .C(_1404_), .Y(_645_) );
NOR2X1 NOR2X1_211 ( .A(_644_), .B(_645_), .Y(_646_) );
INVX1 INVX1_154 ( .A(_142_), .Y(_647_) );
NOR2X1 NOR2X1_212 ( .A(new_wire_586), .B(_647_), .Y(_648_) );
NAND3X1 NAND3X1_158 ( .A(_646_), .B(_648_), .C(_643_), .Y(_649_) );
AOI21X1 AOI21X1_92 ( .A(_630_), .B(_640_), .C(_649_), .Y(_650_) );
NOR2X1 NOR2X1_213 ( .A(new_wire_190), .B(_650_), .Y(_651_) );
OAI21X1 OAI21X1_315 ( .A(_619_), .B(_592_), .C(new_wire_146), .Y(_652_) );
OAI21X1 OAI21X1_316 ( .A(_614_), .B(new_wire_146), .C(_652_), .Y(_1__0_) );
AOI21X1 AOI21X1_93 ( .A(_180_), .B(_185_), .C(new_wire_578), .Y(_653_) );
INVX1 INVX1_155 ( .A(ABL_1_), .Y(_654_) );
AOI22X1 AOI22X1_44 ( .A(new_wire_346), .B(new_wire_92), .C(new_wire_373), .D(new_wire_588), .Y(_655_) );
OAI21X1 OAI21X1_317 ( .A(_654_), .B(new_wire_595), .C(_655_), .Y(_656_) );
AOI21X1 AOI21X1_94 ( .A(new_wire_583), .B(new_wire_346), .C(_656_), .Y(_657_) );
OAI21X1 OAI21X1_318 ( .A(new_wire_349), .B(new_wire_591), .C(_657_), .Y(_658_) );
OR2X2 OR2X2_29 ( .A(_658_), .B(_653_), .Y(_1439__1_) );
OAI21X1 OAI21X1_319 ( .A(_658_), .B(_653_), .C(new_wire_142), .Y(_659_) );
OAI21X1 OAI21X1_320 ( .A(_654_), .B(new_wire_142), .C(_659_), .Y(_1__1_) );
AOI21X1 AOI21X1_95 ( .A(_193_), .B(_198_), .C(new_wire_578), .Y(_660_) );
AOI22X1 AOI22X1_45 ( .A(new_wire_358), .B(new_wire_88), .C(new_wire_368), .D(new_wire_589), .Y(_661_) );
OAI21X1 OAI21X1_321 ( .A(_958_), .B(new_wire_595), .C(_661_), .Y(_662_) );
AOI21X1 AOI21X1_96 ( .A(new_wire_583), .B(new_wire_358), .C(_662_), .Y(_663_) );
OAI21X1 OAI21X1_322 ( .A(new_wire_360), .B(new_wire_591), .C(_663_), .Y(_664_) );
OR2X2 OR2X2_30 ( .A(_664_), .B(_660_), .Y(_1439__2_) );
OAI21X1 OAI21X1_323 ( .A(_664_), .B(_660_), .C(new_wire_150), .Y(_665_) );
OAI21X1 OAI21X1_324 ( .A(_958_), .B(new_wire_150), .C(_665_), .Y(_1__2_) );
AOI21X1 AOI21X1_97 ( .A(_206_), .B(_211_), .C(new_wire_579), .Y(_666_) );
AOI22X1 AOI22X1_46 ( .A(new_wire_352), .B(new_wire_88), .C(new_wire_363), .D(new_wire_589), .Y(_667_) );
OAI21X1 OAI21X1_325 ( .A(_946_), .B(new_wire_595), .C(_667_), .Y(_668_) );
AOI21X1 AOI21X1_98 ( .A(new_wire_584), .B(new_wire_353), .C(_668_), .Y(_669_) );
OAI21X1 OAI21X1_326 ( .A(new_wire_354), .B(new_wire_591), .C(_669_), .Y(_670_) );
OR2X2 OR2X2_31 ( .A(_670_), .B(_666_), .Y(_1439__3_) );
OAI21X1 OAI21X1_327 ( .A(_670_), .B(_666_), .C(new_wire_150), .Y(_671_) );
OAI21X1 OAI21X1_328 ( .A(_946_), .B(new_wire_150), .C(_671_), .Y(_1__3_) );
AOI21X1 AOI21X1_99 ( .A(_219_), .B(_224_), .C(new_wire_579), .Y(_672_) );
AOI22X1 AOI22X1_47 ( .A(new_wire_313), .B(new_wire_92), .C(DIMUX_4_), .D(new_wire_589), .Y(_673_) );
OAI21X1 OAI21X1_329 ( .A(_874_), .B(new_wire_596), .C(_673_), .Y(_674_) );
AOI21X1 AOI21X1_100 ( .A(new_wire_584), .B(new_wire_313), .C(_674_), .Y(_675_) );
OAI21X1 OAI21X1_330 ( .A(new_wire_318), .B(new_wire_592), .C(_675_), .Y(_676_) );
OR2X2 OR2X2_32 ( .A(_676_), .B(_672_), .Y(_1439__4_) );
OAI21X1 OAI21X1_331 ( .A(_676_), .B(_672_), .C(new_wire_148), .Y(_677_) );
OAI21X1 OAI21X1_332 ( .A(_874_), .B(new_wire_148), .C(_677_), .Y(_1__4_) );
AOI21X1 AOI21X1_101 ( .A(_233_), .B(_238_), .C(new_wire_579), .Y(_678_) );
AOI22X1 AOI22X1_48 ( .A(new_wire_296), .B(new_wire_93), .C(new_wire_294), .D(new_wire_589), .Y(_679_) );
OAI21X1 OAI21X1_333 ( .A(_862_), .B(new_wire_596), .C(_679_), .Y(_680_) );
AOI21X1 AOI21X1_102 ( .A(new_wire_584), .B(new_wire_296), .C(_680_), .Y(_681_) );
OAI21X1 OAI21X1_334 ( .A(new_wire_307), .B(new_wire_592), .C(_681_), .Y(_682_) );
OR2X2 OR2X2_33 ( .A(_682_), .B(_678_), .Y(_1439__5_) );
OAI21X1 OAI21X1_335 ( .A(_682_), .B(_678_), .C(new_wire_148), .Y(_683_) );
OAI21X1 OAI21X1_336 ( .A(_862_), .B(new_wire_146), .C(_683_), .Y(_1__5_) );
AOI21X1 AOI21X1_103 ( .A(_246_), .B(_251_), .C(new_wire_579), .Y(_684_) );
AOI22X1 AOI22X1_49 ( .A(new_wire_327), .B(new_wire_90), .C(new_wire_385), .D(new_wire_590), .Y(_685_) );
OAI21X1 OAI21X1_337 ( .A(_895_), .B(new_wire_596), .C(_685_), .Y(_686_) );
AOI21X1 AOI21X1_104 ( .A(new_wire_584), .B(new_wire_327), .C(_686_), .Y(_687_) );
OAI21X1 OAI21X1_338 ( .A(new_wire_328), .B(new_wire_592), .C(_687_), .Y(_688_) );
OR2X2 OR2X2_34 ( .A(_688_), .B(_684_), .Y(_1439__6_) );
OAI21X1 OAI21X1_339 ( .A(_688_), .B(_684_), .C(new_wire_151), .Y(_689_) );
OAI21X1 OAI21X1_340 ( .A(_895_), .B(new_wire_151), .C(_689_), .Y(_1__6_) );
AOI21X1 AOI21X1_105 ( .A(_259_), .B(_264_), .C(new_wire_580), .Y(_690_) );
AOI22X1 AOI22X1_50 ( .A(new_wire_321), .B(new_wire_90), .C(new_wire_388), .D(new_wire_590), .Y(_691_) );
OAI21X1 OAI21X1_341 ( .A(_885_), .B(new_wire_596), .C(_691_), .Y(_692_) );
AOI21X1 AOI21X1_106 ( .A(new_wire_585), .B(new_wire_321), .C(_692_), .Y(_693_) );
OAI21X1 OAI21X1_342 ( .A(new_wire_323), .B(new_wire_592), .C(_693_), .Y(_694_) );
OR2X2 OR2X2_35 ( .A(_694_), .B(_690_), .Y(_1439__7_) );
OAI21X1 OAI21X1_343 ( .A(_694_), .B(_690_), .C(new_wire_148), .Y(_695_) );
OAI21X1 OAI21X1_344 ( .A(_885_), .B(new_wire_146), .C(_695_), .Y(_1__7_) );
OAI21X1 OAI21X1_345 ( .A(_88_), .B(new_wire_538), .C(ABH_0_), .Y(_696_) );
AOI21X1 AOI21X1_107 ( .A(_608_), .B(new_wire_332), .C(_120_), .Y(_697_) );
NAND3X1 NAND3X1_159 ( .A(_696_), .B(_697_), .C(new_wire_580), .Y(_698_) );
OAI21X1 OAI21X1_346 ( .A(_104_), .B(new_wire_581), .C(_595_), .Y(_699_) );
NOR2X1 NOR2X1_214 ( .A(_698_), .B(_699_), .Y(_700_) );
OAI21X1 OAI21X1_347 ( .A(_1008_), .B(new_wire_593), .C(_700_), .Y(_1439__8_) );
NAND2X1 NAND2X1_197 ( .A(_1439__8_), .B(new_wire_142), .Y(_701_) );
OAI21X1 OAI21X1_348 ( .A(_1006_), .B(new_wire_142), .C(_701_), .Y(_0__0_) );
INVX2 INVX2_44 ( .A(new_wire_581), .Y(_702_) );
INVX4 INVX4_7 ( .A(_608_), .Y(_703_) );
OAI21X1 OAI21X1_349 ( .A(new_wire_88), .B(new_wire_586), .C(ABH_1_), .Y(_704_) );
OAI21X1 OAI21X1_350 ( .A(new_wire_348), .B(new_wire_599), .C(_704_), .Y(_705_) );
AOI21X1 AOI21X1_108 ( .A(new_wire_597), .B(new_wire_373), .C(_705_), .Y(_706_) );
OAI21X1 OAI21X1_351 ( .A(_996_), .B(new_wire_593), .C(_706_), .Y(_1439__9_) );
NAND2X1 NAND2X1_198 ( .A(_1439__9_), .B(new_wire_147), .Y(_707_) );
OAI21X1 OAI21X1_352 ( .A(_994_), .B(new_wire_147), .C(_707_), .Y(_0__1_) );
OAI21X1 OAI21X1_353 ( .A(new_wire_89), .B(new_wire_587), .C(ABH_2_), .Y(_708_) );
OAI21X1 OAI21X1_354 ( .A(_360_), .B(new_wire_599), .C(_708_), .Y(_709_) );
AOI21X1 AOI21X1_109 ( .A(new_wire_597), .B(new_wire_369), .C(_709_), .Y(_710_) );
OAI21X1 OAI21X1_355 ( .A(new_wire_370), .B(new_wire_593), .C(_710_), .Y(_1439__10_) );
NAND2X1 NAND2X1_199 ( .A(_1439__10_), .B(new_wire_149), .Y(_711_) );
OAI21X1 OAI21X1_356 ( .A(_981_), .B(new_wire_149), .C(_711_), .Y(_0__2_) );
OAI21X1 OAI21X1_357 ( .A(new_wire_89), .B(new_wire_587), .C(ABH_3_), .Y(_712_) );
OAI21X1 OAI21X1_358 ( .A(_363_), .B(new_wire_599), .C(_712_), .Y(_713_) );
AOI21X1 AOI21X1_110 ( .A(new_wire_597), .B(new_wire_363), .C(_713_), .Y(_714_) );
OAI21X1 OAI21X1_359 ( .A(new_wire_364), .B(new_wire_593), .C(_714_), .Y(_1439__11_) );
NAND2X1 NAND2X1_200 ( .A(_1439__11_), .B(new_wire_143), .Y(_715_) );
OAI21X1 OAI21X1_360 ( .A(_970_), .B(new_wire_143), .C(_715_), .Y(_0__3_) );
OAI22X1 OAI22X1_43 ( .A(_367_), .B(new_wire_599), .C(new_wire_379), .D(new_wire_581), .Y(_716_) );
AOI21X1 AOI21X1_111 ( .A(ABH_4_), .B(_606_), .C(_716_), .Y(_717_) );
OAI21X1 OAI21X1_361 ( .A(new_wire_376), .B(new_wire_594), .C(_717_), .Y(_1439__12_) );
NAND2X1 NAND2X1_201 ( .A(_1439__12_), .B(new_wire_143), .Y(_718_) );
OAI21X1 OAI21X1_362 ( .A(_1020_), .B(new_wire_144), .C(_718_), .Y(_0__4_) );
OAI21X1 OAI21X1_363 ( .A(new_wire_91), .B(new_wire_587), .C(ABH_5_), .Y(_719_) );
OAI21X1 OAI21X1_364 ( .A(new_wire_299), .B(new_wire_600), .C(_719_), .Y(_720_) );
AOI21X1 AOI21X1_112 ( .A(new_wire_597), .B(new_wire_294), .C(_720_), .Y(_721_) );
OAI21X1 OAI21X1_365 ( .A(_787_), .B(new_wire_594), .C(_721_), .Y(_1439__13_) );
NAND2X1 NAND2X1_202 ( .A(_1439__13_), .B(new_wire_144), .Y(_722_) );
OAI21X1 OAI21X1_366 ( .A(_226_), .B(new_wire_144), .C(_722_), .Y(_0__5_) );
INVX1 INVX1_156 ( .A(PC_14_), .Y(_723_) );
OAI21X1 OAI21X1_367 ( .A(new_wire_87), .B(new_wire_587), .C(ABH_6_), .Y(_724_) );
OAI21X1 OAI21X1_368 ( .A(_384_), .B(new_wire_600), .C(_724_), .Y(_725_) );
AOI21X1 AOI21X1_113 ( .A(new_wire_598), .B(new_wire_385), .C(_725_), .Y(_726_) );
OAI21X1 OAI21X1_369 ( .A(_723_), .B(new_wire_594), .C(_726_), .Y(_1439__14_) );
NAND2X1 NAND2X1_203 ( .A(_1439__14_), .B(new_wire_144), .Y(_727_) );
OAI21X1 OAI21X1_370 ( .A(_1049_), .B(new_wire_145), .C(_727_), .Y(_0__6_) );
OAI22X1 OAI22X1_44 ( .A(_387_), .B(new_wire_600), .C(new_wire_387), .D(new_wire_582), .Y(_728_) );
AOI21X1 AOI21X1_114 ( .A(ABH_7_), .B(_606_), .C(_728_), .Y(_729_) );
OAI21X1 OAI21X1_371 ( .A(_1059_), .B(new_wire_594), .C(_729_), .Y(_1439__15_) );
NAND2X1 NAND2X1_204 ( .A(_1439__15_), .B(new_wire_145), .Y(_730_) );
OAI21X1 OAI21X1_372 ( .A(_1061_), .B(new_wire_145), .C(_730_), .Y(_0__7_) );
OAI21X1 OAI21X1_373 ( .A(new_wire_334), .B(new_wire_276), .C(_910_), .Y(_731_) );
NAND2X1 NAND2X1_205 ( .A(_918_), .B(_927_), .Y(_732_) );
NOR2X1 NOR2X1_215 ( .A(_732_), .B(_731_), .Y(_733_) );
INVX1 INVX1_157 ( .A(_902_), .Y(_734_) );
OAI21X1 OAI21X1_374 ( .A(_904_), .B(new_wire_264), .C(_909_), .Y(_735_) );
OAI21X1 OAI21X1_375 ( .A(_735_), .B(_734_), .C(_732_), .Y(_736_) );
NAND2X1 NAND2X1_206 ( .A(new_wire_5), .B(_736_), .Y(_737_) );
OAI22X1 OAI22X1_45 ( .A(new_wire_6), .B(new_wire_334), .C(_733_), .D(_737_), .Y(_9__0_) );
NOR2X1 NOR2X1_216 ( .A(_940_), .B(_928_), .Y(_738_) );
NAND2X1 NAND2X1_207 ( .A(new_wire_16), .B(_1031_), .Y(_739_) );
OAI22X1 OAI22X1_46 ( .A(new_wire_16), .B(new_wire_350), .C(_738_), .D(_739_), .Y(_9__1_) );
INVX1 INVX1_158 ( .A(_1031_), .Y(_740_) );
OAI21X1 OAI21X1_376 ( .A(new_wire_361), .B(new_wire_276), .C(_962_), .Y(_741_) );
NOR2X1 NOR2X1_217 ( .A(_741_), .B(_740_), .Y(_742_) );
NAND3X1 NAND3X1_160 ( .A(_940_), .B(_741_), .C(_928_), .Y(_743_) );
NAND2X1 NAND2X1_208 ( .A(new_wire_17), .B(new_wire_601), .Y(_744_) );
OAI22X1 OAI22X1_47 ( .A(new_wire_7), .B(new_wire_361), .C(_744_), .D(_742_), .Y(_9__2_) );
NOR2X1 NOR2X1_218 ( .A(_1035_), .B(_1032_), .Y(_745_) );
AND2X2 AND2X2_46 ( .A(new_wire_601), .B(_745_), .Y(_746_) );
OAI21X1 OAI21X1_377 ( .A(_745_), .B(new_wire_601), .C(new_wire_17), .Y(_747_) );
OAI22X1 OAI22X1_48 ( .A(new_wire_17), .B(new_wire_355), .C(_746_), .D(_747_), .Y(_9__3_) );
OAI21X1 OAI21X1_378 ( .A(new_wire_319), .B(new_wire_277), .C(_878_), .Y(_748_) );
NOR2X1 NOR2X1_219 ( .A(_745_), .B(new_wire_601), .Y(_749_) );
AOI21X1 AOI21X1_115 ( .A(_749_), .B(_748_), .C(new_wire_186), .Y(_750_) );
OAI21X1 OAI21X1_379 ( .A(_748_), .B(_749_), .C(_750_), .Y(_751_) );
OAI21X1 OAI21X1_380 ( .A(new_wire_7), .B(new_wire_319), .C(_751_), .Y(_9__4_) );
OAI21X1 OAI21X1_381 ( .A(new_wire_307), .B(new_wire_277), .C(_867_), .Y(_752_) );
AOI21X1 AOI21X1_116 ( .A(_749_), .B(_748_), .C(_752_), .Y(_753_) );
INVX1 INVX1_159 ( .A(_879_), .Y(_754_) );
NOR3X1 NOR3X1_15 ( .A(_745_), .B(_754_), .C(new_wire_602), .Y(_755_) );
OR2X2 OR2X2_36 ( .A(new_wire_603), .B(new_wire_186), .Y(_756_) );
OAI22X1 OAI22X1_49 ( .A(new_wire_17), .B(new_wire_308), .C(_753_), .D(_756_), .Y(_9__5_) );
OAI21X1 OAI21X1_382 ( .A(new_wire_328), .B(new_wire_277), .C(_899_), .Y(_757_) );
AOI21X1 AOI21X1_117 ( .A(new_wire_603), .B(_757_), .C(new_wire_186), .Y(_758_) );
OAI21X1 OAI21X1_383 ( .A(_757_), .B(new_wire_603), .C(_758_), .Y(_759_) );
OAI21X1 OAI21X1_384 ( .A(new_wire_18), .B(new_wire_329), .C(_759_), .Y(_9__6_) );
OAI21X1 OAI21X1_385 ( .A(new_wire_323), .B(new_wire_277), .C(_889_), .Y(_760_) );
AOI21X1 AOI21X1_118 ( .A(new_wire_603), .B(_757_), .C(_760_), .Y(_761_) );
NAND3X1 NAND3X1_161 ( .A(_760_), .B(_757_), .C(new_wire_604), .Y(_762_) );
NAND2X1 NAND2X1_209 ( .A(new_wire_6), .B(_762_), .Y(_763_) );
OAI22X1 OAI22X1_50 ( .A(new_wire_6), .B(new_wire_324), .C(_761_), .D(_763_), .Y(_9__7_) );
OAI21X1 OAI21X1_386 ( .A(_1008_), .B(new_wire_278), .C(_1012_), .Y(_764_) );
OAI21X1 OAI21X1_387 ( .A(_901_), .B(_964_), .C(_764_), .Y(_765_) );
NAND3X1 NAND3X1_162 ( .A(_963_), .B(_1030_), .C(_740_), .Y(_766_) );
OR2X2 OR2X2_37 ( .A(_766_), .B(_764_), .Y(_767_) );
NAND3X1 NAND3X1_163 ( .A(new_wire_8), .B(_765_), .C(_767_), .Y(_768_) );
NAND2X1 NAND2X1_210 ( .A(new_wire_186), .B(_1008_), .Y(_769_) );
AND2X2 AND2X2_47 ( .A(_768_), .B(_769_), .Y(_9__8_) );
OAI21X1 OAI21X1_388 ( .A(_996_), .B(new_wire_278), .C(_1000_), .Y(_770_) );
NOR2X1 NOR2X1_220 ( .A(_901_), .B(_964_), .Y(_771_) );
AOI21X1 AOI21X1_119 ( .A(_771_), .B(_764_), .C(_770_), .Y(_772_) );
INVX1 INVX1_160 ( .A(_1013_), .Y(_773_) );
OAI21X1 OAI21X1_389 ( .A(_773_), .B(_766_), .C(new_wire_8), .Y(_774_) );
OAI22X1 OAI22X1_51 ( .A(new_wire_8), .B(_996_), .C(_772_), .D(_774_), .Y(_9__9_) );
OAI21X1 OAI21X1_390 ( .A(new_wire_370), .B(new_wire_278), .C(_987_), .Y(_775_) );
NOR2X1 NOR2X1_221 ( .A(_773_), .B(_766_), .Y(_776_) );
NOR2X1 NOR2X1_222 ( .A(_775_), .B(_776_), .Y(_777_) );
INVX1 INVX1_161 ( .A(_775_), .Y(_778_) );
NAND2X1 NAND2X1_211 ( .A(_1013_), .B(_771_), .Y(_779_) );
OAI21X1 OAI21X1_391 ( .A(_778_), .B(_779_), .C(new_wire_8), .Y(_780_) );
OAI22X1 OAI22X1_52 ( .A(new_wire_9), .B(new_wire_371), .C(_780_), .D(_777_), .Y(_9__10_) );
OAI21X1 OAI21X1_392 ( .A(new_wire_364), .B(new_wire_278), .C(_976_), .Y(_781_) );
AOI21X1 AOI21X1_120 ( .A(_776_), .B(_775_), .C(_781_), .Y(_782_) );
OAI21X1 OAI21X1_393 ( .A(_1014_), .B(_766_), .C(new_wire_9), .Y(_783_) );
OAI22X1 OAI22X1_53 ( .A(new_wire_9), .B(new_wire_365), .C(_783_), .D(_782_), .Y(_9__11_) );
NOR2X1 NOR2X1_223 ( .A(new_wire_380), .B(_1015_), .Y(_784_) );
INVX1 INVX1_162 ( .A(new_wire_381), .Y(_785_) );
OAI21X1 OAI21X1_394 ( .A(_785_), .B(_1043_), .C(new_wire_18), .Y(_786_) );
OAI22X1 OAI22X1_54 ( .A(new_wire_18), .B(new_wire_377), .C(_784_), .D(_786_), .Y(_9__12_) );
BUFX2 BUFX2_17 ( .A(_1439__0_), .Y(AB[0]) );
BUFX2 BUFX2_18 ( .A(_1439__1_), .Y(AB[1]) );
BUFX2 BUFX2_19 ( .A(_1439__2_), .Y(AB[2]) );
BUFX2 BUFX2_20 ( .A(_1439__3_), .Y(AB[3]) );
BUFX2 BUFX2_21 ( .A(_1439__4_), .Y(AB[4]) );
BUFX2 BUFX2_22 ( .A(_1439__5_), .Y(AB[5]) );
BUFX2 BUFX2_23 ( .A(_1439__6_), .Y(AB[6]) );
BUFX2 BUFX2_24 ( .A(_1439__7_), .Y(AB[7]) );
BUFX2 BUFX2_25 ( .A(_1439__8_), .Y(AB[8]) );
BUFX2 BUFX2_26 ( .A(_1439__9_), .Y(AB[9]) );
BUFX2 BUFX2_27 ( .A(_1439__10_), .Y(AB[10]) );
BUFX2 BUFX2_28 ( .A(_1439__11_), .Y(AB[11]) );
BUFX2 BUFX2_29 ( .A(_1439__12_), .Y(AB[12]) );
BUFX2 BUFX2_30 ( .A(_1439__13_), .Y(AB[13]) );
BUFX2 BUFX2_31 ( .A(_1439__14_), .Y(AB[14]) );
BUFX2 BUFX2_32 ( .A(_1439__15_), .Y(AB[15]) );
BUFX2 BUFX2_33 ( .A(_1440__0_), .Y(DO[0]) );
BUFX2 BUFX2_34 ( .A(_1440__1_), .Y(DO[1]) );
BUFX2 BUFX2_35 ( .A(_1440__2_), .Y(DO[2]) );
BUFX2 BUFX2_36 ( .A(_1440__3_), .Y(DO[3]) );
BUFX2 BUFX2_37 ( .A(_1440__4_), .Y(DO[4]) );
BUFX2 BUFX2_38 ( .A(_1440__5_), .Y(DO[5]) );
BUFX2 BUFX2_39 ( .A(_1440__6_), .Y(DO[6]) );
BUFX2 BUFX2_40 ( .A(_1440__7_), .Y(DO[7]) );
BUFX2 BUFX2_41 ( .A(_1441_), .Y(WE) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(new_wire_49), .D(_1443__0_), .Q(AXYS_0__0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(new_wire_58), .D(_1443__1_), .Q(AXYS_0__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(new_wire_40), .D(_1443__2_), .Q(AXYS_0__2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(new_wire_52), .D(_1443__3_), .Q(AXYS_0__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(new_wire_58), .D(_1443__4_), .Q(AXYS_0__4_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(new_wire_49), .D(_1443__5_), .Q(AXYS_0__5_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(new_wire_49), .D(_1443__6_), .Q(AXYS_0__6_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(new_wire_40), .D(_1443__7_), .Q(AXYS_0__7_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(new_wire_58), .D(_1442__0_), .Q(AXYS_1__0_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(new_wire_52), .D(_1442__1_), .Q(AXYS_1__1_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(new_wire_40), .D(_1442__2_), .Q(AXYS_1__2_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(new_wire_49), .D(_1442__3_), .Q(AXYS_1__3_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(new_wire_58), .D(_1442__4_), .Q(AXYS_1__4_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(new_wire_50), .D(_1442__5_), .Q(AXYS_1__5_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(new_wire_50), .D(_1442__6_), .Q(AXYS_1__6_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(new_wire_40), .D(_1442__7_), .Q(AXYS_1__7_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(new_wire_50), .D(_1445__0_), .Q(AXYS_3__0_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(new_wire_59), .D(_1445__1_), .Q(AXYS_3__1_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(new_wire_41), .D(_1445__2_), .Q(AXYS_3__2_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(new_wire_41), .D(_1445__3_), .Q(AXYS_3__3_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(new_wire_59), .D(_1445__4_), .Q(AXYS_3__4_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(new_wire_41), .D(_1445__5_), .Q(AXYS_3__5_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(new_wire_50), .D(_1445__6_), .Q(AXYS_3__6_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(new_wire_41), .D(_1445__7_), .Q(AXYS_3__7_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(new_wire_51), .D(_1444__0_), .Q(AXYS_2__0_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(new_wire_59), .D(_1444__1_), .Q(AXYS_2__1_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(new_wire_42), .D(_1444__2_), .Q(AXYS_2__2_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(new_wire_55), .D(_1444__3_), .Q(AXYS_2__3_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(new_wire_59), .D(_1444__4_), .Q(AXYS_2__4_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(new_wire_60), .D(_1444__5_), .Q(AXYS_2__5_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(new_wire_51), .D(_1444__6_), .Q(AXYS_2__6_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(new_wire_42), .D(_1444__7_), .Q(AXYS_2__7_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(new_wire_52), .D(_7_), .Q(NMI_edge) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(new_wire_42), .D(NMI), .Q(NMI_1) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(new_wire_43), .D(_22__0_), .Q(cond_code_0_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(new_wire_43), .D(_22__1_), .Q(cond_code_1_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(new_wire_46), .D(_22__2_), .Q(cond_code_2_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(new_wire_43), .D(_30_), .Q(plp) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(new_wire_43), .D(_29_), .Q(php) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(new_wire_70), .D(_17_), .Q(clc) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(new_wire_64), .D(_33_), .Q(sec) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(new_wire_70), .D(_18_), .Q(cld) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(new_wire_70), .D(_34_), .Q(sed) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(new_wire_70), .D(_19_), .Q(cli) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(new_wire_71), .D(_35_), .Q(sei) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(new_wire_44), .D(_20_), .Q(clv) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(new_wire_64), .D(_16_), .Q(bit_ins) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(new_wire_64), .D(_28__0_), .Q(op_0_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(new_wire_64), .D(_28__1_), .Q(op_1_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(new_wire_65), .D(_28__2_), .Q(op_2_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(new_wire_65), .D(_28__3_), .Q(op_3_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(new_wire_71), .D(_32_), .Q(rotate) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(new_wire_65), .D(_37_), .Q(shift_right) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(new_wire_71), .D(_21_), .Q(compare) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(new_wire_44), .D(_36_), .Q(shift) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(new_wire_55), .D(_12_), .Q(adc_bcd) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(new_wire_55), .D(_13_), .Q(adc_sbc) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(new_wire_71), .D(_24_), .Q(inc) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(new_wire_65), .D(_26_), .Q(load_only) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(new_wire_44), .D(_40_), .Q(write_back) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(new_wire_44), .D(_39_), .Q(store) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(new_wire_45), .D(_25_), .Q(index_y) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(new_wire_45), .D(_38__0_), .Q(src_reg_0_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(new_wire_72), .D(_38__1_), .Q(src_reg_1_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(new_wire_46), .D(_23__0_), .Q(dst_reg_0_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(new_wire_45), .D(_23__1_), .Q(dst_reg_1_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(new_wire_45), .D(_27_), .Q(load_reg) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(new_wire_61), .D(_31_), .Q(res) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(new_wire_67), .D(new_wire_375), .Q(DIHOLD_0_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(new_wire_61), .D(new_wire_373), .Q(DIHOLD_1_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(new_wire_52), .D(new_wire_369), .Q(DIHOLD_2_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(new_wire_67), .D(new_wire_363), .Q(DIHOLD_3_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(new_wire_53), .D(DIMUX_4_), .Q(DIHOLD_4_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(new_wire_67), .D(new_wire_294), .Q(DIHOLD_5_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(new_wire_46), .D(new_wire_385), .Q(DIHOLD_6_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(new_wire_46), .D(new_wire_389), .Q(DIHOLD_7_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(new_wire_55), .D(_4__0_), .Q(IRHOLD_0_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(new_wire_56), .D(_4__1_), .Q(IRHOLD_1_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(new_wire_47), .D(_4__2_), .Q(IRHOLD_2_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(new_wire_56), .D(_4__3_), .Q(IRHOLD_3_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(new_wire_56), .D(_4__4_), .Q(IRHOLD_4_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(new_wire_56), .D(_4__5_), .Q(IRHOLD_5_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(new_wire_47), .D(_4__6_), .Q(IRHOLD_6_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(new_wire_72), .D(_4__7_), .Q(IRHOLD_7_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(new_wire_57), .D(_5_), .Q(IRHOLD_valid) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(new_wire_47), .D(_10_), .Q(V) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(new_wire_47), .D(_3_), .Q(D) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(new_wire_53), .D(_6_), .Q(I) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(new_wire_48), .D(_8_), .Q(N) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(new_wire_48), .D(_11_), .Q(Z) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(new_wire_48), .D(_2_), .Q(C) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(new_wire_48), .D(_15_), .Q(backwards) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(new_wire_57), .D(_14_), .Q(adj_bcd) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(new_wire_67), .D(_1__0_), .Q(ABL_0_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(new_wire_73), .D(_1__1_), .Q(ABL_1_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(new_wire_68), .D(_1__2_), .Q(ABL_2_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(new_wire_68), .D(_1__3_), .Q(ABL_3_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(new_wire_68), .D(_1__4_), .Q(ABL_4_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(new_wire_68), .D(_1__5_), .Q(ABL_5_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(new_wire_42), .D(_1__6_), .Q(ABL_6_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(new_wire_69), .D(_1__7_), .Q(ABL_7_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(new_wire_53), .D(_0__0_), .Q(ABH_0_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(new_wire_73), .D(_0__1_), .Q(ABH_1_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(new_wire_69), .D(_0__2_), .Q(ABH_2_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(new_wire_53), .D(_0__3_), .Q(ABH_3_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(new_wire_54), .D(_0__4_), .Q(ABH_4_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(new_wire_54), .D(_0__5_), .Q(ABH_5_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(new_wire_54), .D(_0__6_), .Q(ABH_6_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(new_wire_54), .D(_0__7_), .Q(ABH_7_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(new_wire_61), .D(_9__0_), .Q(PC_0_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(new_wire_73), .D(_9__1_), .Q(PC_1_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(new_wire_73), .D(_9__2_), .Q(PC_2_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(new_wire_74), .D(_9__3_), .Q(PC_3_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(new_wire_69), .D(_9__4_), .Q(PC_4_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(new_wire_74), .D(_9__5_), .Q(PC_5_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(new_wire_61), .D(_9__6_), .Q(PC_6_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(new_wire_62), .D(_9__7_), .Q(PC_7_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(new_wire_74), .D(_9__8_), .Q(PC_8_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(new_wire_74), .D(_9__9_), .Q(PC_9_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(new_wire_75), .D(_9__10_), .Q(PC_10_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(new_wire_69), .D(_9__11_), .Q(PC_11_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(new_wire_75), .D(_9__12_), .Q(PC_12_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(new_wire_75), .D(_9__13_), .Q(PC_13_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(new_wire_62), .D(_9__14_), .Q(PC_14_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(new_wire_75), .D(_9__15_), .Q(PC_15_) );
DFFSR DFFSR_1 ( .CLK(new_wire_62), .D(_1438__0_), .Q(state_0_), .R(new_wire_545), .S(vdd) );
DFFSR DFFSR_2 ( .CLK(new_wire_62), .D(_1438__1_), .Q(state_1_), .R(new_wire_545), .S(vdd) );
DFFSR DFFSR_3 ( .CLK(new_wire_63), .D(_1438__2_), .Q(state_2_), .R(new_wire_545), .S(vdd) );
DFFSR DFFSR_4 ( .CLK(new_wire_63), .D(_1438__3_), .Q(state_3_), .R(vdd), .S(new_wire_546) );
DFFSR DFFSR_5 ( .CLK(new_wire_63), .D(_1438__4_), .Q(state_4_), .R(new_wire_546), .S(vdd) );
DFFSR DFFSR_6 ( .CLK(new_wire_63), .D(_1438__5_), .Q(state_5_), .R(new_wire_546), .S(vdd) );
OR2X2 OR2X2_38 ( .A(new_wire_353), .B(new_wire_332), .Y(_1626_) );
NOR2X1 NOR2X1_224 ( .A(new_wire_327), .B(new_wire_322), .Y(_1627_) );
NOR2X1 NOR2X1_225 ( .A(new_wire_314), .B(new_wire_296), .Y(_1628_) );
NOR2X1 NOR2X1_226 ( .A(new_wire_358), .B(new_wire_346), .Y(_1629_) );
NAND3X1 NAND3X1_164 ( .A(_1627_), .B(_1628_), .C(_1629_), .Y(_1630_) );
NOR2X1 NOR2X1_227 ( .A(_1626_), .B(_1630_), .Y(AZ) );
INVX8 INVX8_7 ( .A(new_wire_12), .Y(_1631_) );
NAND2X1 NAND2X1_212 ( .A(new_wire_336), .B(new_wire_166), .Y(_1632_) );
INVX2 INVX2_45 ( .A(new_wire_531), .Y(_1633_) );
NOR2X1 NOR2X1_228 ( .A(new_wire_527), .B(new_wire_605), .Y(_1634_) );
INVX1 INVX1_163 ( .A(new_wire_524), .Y(_1635_) );
NOR2X1 NOR2X1_229 ( .A(alu_op_1_), .B(_1635_), .Y(_1636_) );
INVX1 INVX1_164 ( .A(BI_5_), .Y(_1637_) );
NOR2X1 NOR2X1_230 ( .A(new_wire_524), .B(_1637_), .Y(_1638_) );
INVX4 INVX4_8 ( .A(alu_op_1_), .Y(_1639_) );
INVX1 INVX1_165 ( .A(AI_5_), .Y(_1640_) );
OAI21X1 OAI21X1_395 ( .A(new_wire_610), .B(_1640_), .C(BI_5_), .Y(_1641_) );
OAI21X1 OAI21X1_396 ( .A(_1636_), .B(_1638_), .C(_1641_), .Y(_1642_) );
INVX1 INVX1_166 ( .A(_1638_), .Y(_1643_) );
AOI21X1 AOI21X1_121 ( .A(_1643_), .B(_1640_), .C(new_wire_553), .Y(_1644_) );
AOI22X1 AOI22X1_51 ( .A(new_wire_553), .B(AI_6_), .C(_1642_), .D(_1644_), .Y(_1645_) );
INVX1 INVX1_167 ( .A(_1645_), .Y(_1646_) );
INVX1 INVX1_168 ( .A(new_wire_527), .Y(_1647_) );
NOR2X1 NOR2X1_231 ( .A(new_wire_531), .B(_1647_), .Y(_1648_) );
OAI21X1 OAI21X1_397 ( .A(new_wire_527), .B(new_wire_531), .C(BI_5_), .Y(_1649_) );
OAI21X1 OAI21X1_398 ( .A(BI_5_), .B(new_wire_612), .C(_1649_), .Y(_1650_) );
INVX1 INVX1_169 ( .A(_1650_), .Y(_1651_) );
OAI21X1 OAI21X1_399 ( .A(new_wire_607), .B(_1651_), .C(_1646_), .Y(_1652_) );
INVX1 INVX1_170 ( .A(new_wire_614), .Y(_1653_) );
INVX2 INVX2_46 ( .A(new_wire_553), .Y(_1654_) );
NAND2X1 NAND2X1_213 ( .A(new_wire_524), .B(new_wire_610), .Y(_1655_) );
AND2X2 AND2X2_48 ( .A(_1635_), .B(BI_4_), .Y(_1656_) );
NAND2X1 NAND2X1_214 ( .A(AI_4_), .B(_1656_), .Y(_1657_) );
AOI22X1 AOI22X1_52 ( .A(new_wire_610), .B(BI_4_), .C(_1655_), .D(_1657_), .Y(_1658_) );
OAI21X1 OAI21X1_400 ( .A(AI_4_), .B(_1656_), .C(new_wire_616), .Y(_1659_) );
OAI22X1 OAI22X1_55 ( .A(new_wire_616), .B(_1640_), .C(_1659_), .D(_1658_), .Y(_1660_) );
OAI21X1 OAI21X1_401 ( .A(new_wire_527), .B(new_wire_531), .C(BI_4_), .Y(_1661_) );
OAI21X1 OAI21X1_402 ( .A(BI_4_), .B(new_wire_612), .C(_1661_), .Y(_1662_) );
INVX1 INVX1_171 ( .A(_1662_), .Y(_1663_) );
OAI21X1 OAI21X1_403 ( .A(new_wire_607), .B(_1663_), .C(_1660_), .Y(_1664_) );
INVX1 INVX1_172 ( .A(AI_3_), .Y(_1665_) );
INVX1 INVX1_173 ( .A(BI_2_), .Y(_1666_) );
NOR2X1 NOR2X1_232 ( .A(new_wire_524), .B(_1666_), .Y(_1667_) );
INVX1 INVX1_174 ( .A(AI_2_), .Y(_1668_) );
OAI21X1 OAI21X1_404 ( .A(new_wire_610), .B(_1668_), .C(BI_2_), .Y(_1669_) );
OAI21X1 OAI21X1_405 ( .A(_1636_), .B(_1667_), .C(_1669_), .Y(_1670_) );
OAI21X1 OAI21X1_406 ( .A(new_wire_525), .B(_1666_), .C(_1668_), .Y(_1671_) );
NAND3X1 NAND3X1_165 ( .A(new_wire_616), .B(_1671_), .C(_1670_), .Y(_1452_) );
OAI21X1 OAI21X1_407 ( .A(new_wire_616), .B(_1665_), .C(_1452_), .Y(_1453_) );
OAI21X1 OAI21X1_408 ( .A(new_wire_528), .B(new_wire_532), .C(BI_2_), .Y(_1454_) );
OAI21X1 OAI21X1_409 ( .A(BI_2_), .B(new_wire_612), .C(_1454_), .Y(_1455_) );
OAI21X1 OAI21X1_410 ( .A(new_wire_528), .B(new_wire_605), .C(_1455_), .Y(_1456_) );
NAND3X1 NAND3X1_166 ( .A(AI_1_), .B(new_wire_506), .C(_1635_), .Y(_1457_) );
AOI22X1 AOI22X1_53 ( .A(new_wire_611), .B(new_wire_506), .C(_1655_), .D(_1457_), .Y(_1458_) );
INVX1 INVX1_175 ( .A(AI_1_), .Y(_1459_) );
INVX1 INVX1_176 ( .A(new_wire_506), .Y(_1460_) );
OAI21X1 OAI21X1_411 ( .A(new_wire_525), .B(_1460_), .C(_1459_), .Y(_1461_) );
NAND2X1 NAND2X1_215 ( .A(new_wire_617), .B(_1461_), .Y(_1462_) );
OAI22X1 OAI22X1_56 ( .A(new_wire_617), .B(_1668_), .C(_1462_), .D(_1458_), .Y(_1463_) );
OAI21X1 OAI21X1_412 ( .A(new_wire_528), .B(new_wire_532), .C(new_wire_506), .Y(_1464_) );
OAI21X1 OAI21X1_413 ( .A(new_wire_507), .B(new_wire_612), .C(_1464_), .Y(_1465_) );
INVX1 INVX1_177 ( .A(_1465_), .Y(_1466_) );
OAI21X1 OAI21X1_414 ( .A(new_wire_607), .B(_1466_), .C(_1463_), .Y(_1467_) );
NAND2X1 NAND2X1_216 ( .A(new_wire_553), .B(AI_1_), .Y(_1468_) );
NAND2X1 NAND2X1_217 ( .A(new_wire_504), .B(_1635_), .Y(_1469_) );
NAND2X1 NAND2X1_218 ( .A(alu_op_1_), .B(AI_0_), .Y(_1470_) );
AOI22X1 AOI22X1_54 ( .A(new_wire_504), .B(_1470_), .C(_1655_), .D(_1469_), .Y(_1471_) );
INVX1 INVX1_178 ( .A(AI_0_), .Y(_1472_) );
INVX1 INVX1_179 ( .A(new_wire_504), .Y(_1473_) );
OAI21X1 OAI21X1_415 ( .A(new_wire_525), .B(_1473_), .C(_1472_), .Y(_1474_) );
NAND2X1 NAND2X1_219 ( .A(new_wire_617), .B(_1474_), .Y(_1475_) );
OAI21X1 OAI21X1_416 ( .A(_1471_), .B(_1475_), .C(_1468_), .Y(_1476_) );
OAI21X1 OAI21X1_417 ( .A(new_wire_528), .B(new_wire_532), .C(new_wire_504), .Y(_1477_) );
OAI21X1 OAI21X1_418 ( .A(new_wire_505), .B(new_wire_613), .C(_1477_), .Y(_1478_) );
OAI21X1 OAI21X1_419 ( .A(new_wire_529), .B(new_wire_605), .C(_1478_), .Y(_1479_) );
OAI21X1 OAI21X1_420 ( .A(_1647_), .B(new_wire_605), .C(CI), .Y(_1480_) );
NOR2X1 NOR2X1_233 ( .A(new_wire_554), .B(_1480_), .Y(_1481_) );
MUX2X1 MUX2X1_35 ( .A(alu_op_1_), .B(_1473_), .S(new_wire_525), .Y(_1482_) );
NAND2X1 NAND2X1_220 ( .A(new_wire_505), .B(_1470_), .Y(_1483_) );
NAND2X1 NAND2X1_221 ( .A(_1483_), .B(_1482_), .Y(_1484_) );
AOI21X1 AOI21X1_122 ( .A(_1469_), .B(_1472_), .C(new_wire_554), .Y(_1485_) );
NAND2X1 NAND2X1_222 ( .A(_1485_), .B(_1484_), .Y(_1486_) );
NAND3X1 NAND3X1_167 ( .A(_1468_), .B(_1478_), .C(_1486_), .Y(_1487_) );
AOI22X1 AOI22X1_55 ( .A(_1476_), .B(_1479_), .C(_1481_), .D(_1487_), .Y(_1488_) );
NOR2X1 NOR2X1_234 ( .A(_1466_), .B(_1463_), .Y(_1489_) );
OAI21X1 OAI21X1_421 ( .A(_1489_), .B(_1488_), .C(_1467_), .Y(_1490_) );
MUX2X1 MUX2X1_36 ( .A(_1456_), .B(_1455_), .S(_1453_), .Y(_1491_) );
AOI22X1 AOI22X1_56 ( .A(_1453_), .B(_1456_), .C(_1491_), .D(_1490_), .Y(_1492_) );
NAND2X1 NAND2X1_223 ( .A(new_wire_554), .B(AI_4_), .Y(_1493_) );
INVX1 INVX1_180 ( .A(BI_3_), .Y(_1494_) );
NOR2X1 NOR2X1_235 ( .A(new_wire_526), .B(_1494_), .Y(_1495_) );
NAND2X1 NAND2X1_224 ( .A(AI_3_), .B(_1495_), .Y(_1496_) );
AOI22X1 AOI22X1_57 ( .A(new_wire_611), .B(BI_3_), .C(_1655_), .D(_1496_), .Y(_1497_) );
OAI21X1 OAI21X1_422 ( .A(AI_3_), .B(_1495_), .C(new_wire_617), .Y(_1498_) );
OAI21X1 OAI21X1_423 ( .A(_1498_), .B(_1497_), .C(_1493_), .Y(_1499_) );
OAI21X1 OAI21X1_424 ( .A(new_wire_532), .B(_1647_), .C(_1494_), .Y(_1500_) );
OAI21X1 OAI21X1_425 ( .A(new_wire_529), .B(new_wire_533), .C(BI_3_), .Y(_1501_) );
AND2X2 AND2X2_49 ( .A(_1500_), .B(_1501_), .Y(_1502_) );
OAI21X1 OAI21X1_426 ( .A(new_wire_607), .B(_1502_), .C(_1499_), .Y(_1503_) );
OAI21X1 OAI21X1_427 ( .A(_1499_), .B(_1502_), .C(_1503_), .Y(_1504_) );
XOR2X1 XOR2X1_2 ( .A(_1492_), .B(_1504_), .Y(_1505_) );
INVX1 INVX1_181 ( .A(ALU_BCD), .Y(_1506_) );
INVX1 INVX1_182 ( .A(_1478_), .Y(_1507_) );
OAI21X1 OAI21X1_428 ( .A(new_wire_608), .B(_1507_), .C(_1476_), .Y(_1508_) );
INVX1 INVX1_183 ( .A(_1481_), .Y(_1509_) );
NOR2X1 NOR2X1_236 ( .A(_1507_), .B(_1476_), .Y(_1510_) );
OAI21X1 OAI21X1_429 ( .A(_1509_), .B(_1510_), .C(_1508_), .Y(_1511_) );
OAI21X1 OAI21X1_430 ( .A(new_wire_529), .B(new_wire_606), .C(_1465_), .Y(_1512_) );
AOI21X1 AOI21X1_123 ( .A(_1463_), .B(_1512_), .C(_1489_), .Y(_1513_) );
NAND2X1 NAND2X1_225 ( .A(_1513_), .B(_1511_), .Y(_1514_) );
OAI21X1 OAI21X1_431 ( .A(_1463_), .B(_1466_), .C(_1467_), .Y(_1515_) );
NAND2X1 NAND2X1_226 ( .A(_1488_), .B(_1515_), .Y(_1516_) );
NAND2X1 NAND2X1_227 ( .A(_1516_), .B(_1514_), .Y(_1517_) );
NAND2X1 NAND2X1_228 ( .A(_1491_), .B(_1490_), .Y(_1518_) );
INVX1 INVX1_184 ( .A(_1455_), .Y(_1519_) );
OAI21X1 OAI21X1_432 ( .A(new_wire_608), .B(_1519_), .C(_1453_), .Y(_1520_) );
OAI21X1 OAI21X1_433 ( .A(_1453_), .B(_1519_), .C(_1520_), .Y(_1521_) );
NAND3X1 NAND3X1_168 ( .A(_1467_), .B(_1521_), .C(_1514_), .Y(_1522_) );
NAND2X1 NAND2X1_229 ( .A(_1518_), .B(_1522_), .Y(_1523_) );
AOI21X1 AOI21X1_124 ( .A(_1523_), .B(_1517_), .C(_1506_), .Y(_1524_) );
OAI21X1 OAI21X1_434 ( .A(_1504_), .B(_1492_), .C(_1503_), .Y(_1525_) );
AOI21X1 AOI21X1_125 ( .A(_1524_), .B(_1505_), .C(_1525_), .Y(_1526_) );
OAI21X1 OAI21X1_435 ( .A(_1660_), .B(_1663_), .C(_1664_), .Y(_1527_) );
OAI21X1 OAI21X1_436 ( .A(_1527_), .B(_1526_), .C(_1664_), .Y(_1528_) );
OAI21X1 OAI21X1_437 ( .A(_1646_), .B(_1651_), .C(new_wire_614), .Y(_1529_) );
INVX1 INVX1_185 ( .A(_1529_), .Y(_1530_) );
AOI21X1 AOI21X1_126 ( .A(_1528_), .B(_1530_), .C(_1653_), .Y(_1531_) );
INVX1 INVX1_186 ( .A(BI_7_), .Y(_1532_) );
NOR2X1 NOR2X1_237 ( .A(new_wire_526), .B(_1532_), .Y(_1533_) );
INVX1 INVX1_187 ( .A(AI_7_), .Y(_1534_) );
OAI21X1 OAI21X1_438 ( .A(new_wire_611), .B(_1534_), .C(BI_7_), .Y(_1535_) );
OAI21X1 OAI21X1_439 ( .A(_1636_), .B(_1533_), .C(_1535_), .Y(_1536_) );
INVX1 INVX1_188 ( .A(_1533_), .Y(_1537_) );
AOI21X1 AOI21X1_127 ( .A(_1537_), .B(_1534_), .C(new_wire_554), .Y(_1538_) );
AOI22X1 AOI22X1_58 ( .A(CI), .B(new_wire_555), .C(_1536_), .D(_1538_), .Y(_1539_) );
INVX1 INVX1_189 ( .A(_1539_), .Y(_1540_) );
OAI21X1 OAI21X1_440 ( .A(new_wire_529), .B(new_wire_533), .C(BI_7_), .Y(_1541_) );
OAI21X1 OAI21X1_441 ( .A(BI_7_), .B(new_wire_613), .C(_1541_), .Y(_1542_) );
INVX1 INVX1_190 ( .A(_1542_), .Y(_1543_) );
OAI21X1 OAI21X1_442 ( .A(_1543_), .B(new_wire_608), .C(_1540_), .Y(_1544_) );
INVX1 INVX1_191 ( .A(_1544_), .Y(_1545_) );
INVX1 INVX1_192 ( .A(BI_6_), .Y(_1546_) );
NOR2X1 NOR2X1_238 ( .A(new_wire_526), .B(_1546_), .Y(_1547_) );
INVX1 INVX1_193 ( .A(AI_6_), .Y(_1548_) );
OAI21X1 OAI21X1_443 ( .A(new_wire_611), .B(_1548_), .C(BI_6_), .Y(_1549_) );
OAI21X1 OAI21X1_444 ( .A(_1636_), .B(_1547_), .C(_1549_), .Y(_1550_) );
INVX1 INVX1_194 ( .A(_1547_), .Y(_1551_) );
AOI21X1 AOI21X1_128 ( .A(_1551_), .B(_1548_), .C(new_wire_555), .Y(_1552_) );
AOI22X1 AOI22X1_59 ( .A(AI_7_), .B(new_wire_555), .C(_1550_), .D(_1552_), .Y(_1553_) );
INVX1 INVX1_195 ( .A(_1553_), .Y(_1554_) );
OAI21X1 OAI21X1_445 ( .A(new_wire_530), .B(new_wire_533), .C(BI_6_), .Y(_1555_) );
OAI21X1 OAI21X1_446 ( .A(BI_6_), .B(new_wire_613), .C(_1555_), .Y(_1556_) );
INVX1 INVX1_196 ( .A(_1556_), .Y(_1557_) );
OAI21X1 OAI21X1_447 ( .A(new_wire_608), .B(_1557_), .C(_1554_), .Y(_1558_) );
INVX1 INVX1_197 ( .A(_1558_), .Y(_1559_) );
OAI21X1 OAI21X1_448 ( .A(_1540_), .B(_1543_), .C(_1544_), .Y(_1560_) );
INVX1 INVX1_198 ( .A(_1560_), .Y(_1561_) );
AOI21X1 AOI21X1_129 ( .A(_1561_), .B(_1559_), .C(_1545_), .Y(_1562_) );
OAI21X1 OAI21X1_449 ( .A(_1554_), .B(_1557_), .C(_1558_), .Y(_1563_) );
INVX1 INVX1_199 ( .A(_1563_), .Y(_1564_) );
NAND2X1 NAND2X1_230 ( .A(_1564_), .B(_1561_), .Y(_1565_) );
OAI21X1 OAI21X1_450 ( .A(_1565_), .B(_1531_), .C(_1562_), .Y(_1566_) );
NAND3X1 NAND3X1_169 ( .A(new_wire_555), .B(AI_0_), .C(_1566_), .Y(_1567_) );
NAND2X1 NAND2X1_231 ( .A(new_wire_556), .B(AI_0_), .Y(_1568_) );
OR2X2 OR2X2_39 ( .A(_1531_), .B(_1565_), .Y(_1569_) );
NAND3X1 NAND3X1_170 ( .A(_1568_), .B(_1562_), .C(_1569_), .Y(_1570_) );
INVX1 INVX1_200 ( .A(_1664_), .Y(_1571_) );
NAND2X1 NAND2X1_232 ( .A(_1505_), .B(_1524_), .Y(_1572_) );
INVX1 INVX1_201 ( .A(_1525_), .Y(_1573_) );
INVX1 INVX1_202 ( .A(_1660_), .Y(_1574_) );
INVX1 INVX1_203 ( .A(new_wire_609), .Y(_1575_) );
OAI21X1 OAI21X1_451 ( .A(_1575_), .B(_1574_), .C(_1662_), .Y(_1576_) );
OR2X2 OR2X2_40 ( .A(_1576_), .B(_1574_), .Y(_1577_) );
NAND2X1 NAND2X1_233 ( .A(_1574_), .B(_1576_), .Y(_1578_) );
AOI22X1 AOI22X1_60 ( .A(_1577_), .B(_1578_), .C(_1573_), .D(_1572_), .Y(_1579_) );
OAI21X1 OAI21X1_452 ( .A(_1571_), .B(_1579_), .C(_1530_), .Y(_1580_) );
OAI21X1 OAI21X1_453 ( .A(_1575_), .B(_1553_), .C(_1556_), .Y(_1581_) );
OR2X2 OR2X2_41 ( .A(_1581_), .B(_1553_), .Y(_1582_) );
NAND2X1 NAND2X1_234 ( .A(_1553_), .B(_1581_), .Y(_1583_) );
AOI22X1 AOI22X1_61 ( .A(_1582_), .B(_1583_), .C(new_wire_614), .D(_1580_), .Y(_1584_) );
OAI21X1 OAI21X1_454 ( .A(_1559_), .B(_1584_), .C(_1560_), .Y(_1585_) );
OAI21X1 OAI21X1_455 ( .A(new_wire_530), .B(new_wire_606), .C(_1662_), .Y(_1586_) );
XNOR2X1 XNOR2X1_8 ( .A(_1492_), .B(_1504_), .Y(_1587_) );
NAND3X1 NAND3X1_171 ( .A(_1467_), .B(_1491_), .C(_1514_), .Y(_1588_) );
NAND2X1 NAND2X1_235 ( .A(_1521_), .B(_1490_), .Y(_1589_) );
NAND3X1 NAND3X1_172 ( .A(_1589_), .B(_1517_), .C(_1588_), .Y(_1590_) );
NAND2X1 NAND2X1_236 ( .A(ALU_BCD), .B(_1590_), .Y(_1591_) );
OAI21X1 OAI21X1_456 ( .A(_1591_), .B(_1587_), .C(_1573_), .Y(_1592_) );
INVX1 INVX1_204 ( .A(_1527_), .Y(_1593_) );
AOI22X1 AOI22X1_62 ( .A(_1660_), .B(_1586_), .C(_1593_), .D(_1592_), .Y(_1594_) );
OAI21X1 OAI21X1_457 ( .A(_1529_), .B(_1594_), .C(new_wire_614), .Y(_1595_) );
NAND2X1 NAND2X1_237 ( .A(_1564_), .B(_1595_), .Y(_1596_) );
NAND3X1 NAND3X1_173 ( .A(_1558_), .B(_1561_), .C(_1596_), .Y(_1597_) );
NAND2X1 NAND2X1_238 ( .A(_1597_), .B(_1585_), .Y(_1598_) );
NAND2X1 NAND2X1_239 ( .A(_1529_), .B(_1594_), .Y(_1599_) );
NAND2X1 NAND2X1_240 ( .A(_1599_), .B(_1580_), .Y(_1600_) );
NAND3X1 NAND3X1_174 ( .A(new_wire_615), .B(_1563_), .C(_1580_), .Y(_1601_) );
NAND2X1 NAND2X1_241 ( .A(_1601_), .B(_1596_), .Y(_1602_) );
AOI21X1 AOI21X1_130 ( .A(_1602_), .B(_1600_), .C(_1506_), .Y(_1603_) );
AOI22X1 AOI22X1_63 ( .A(_1567_), .B(_1570_), .C(_1598_), .D(_1603_), .Y(_1604_) );
OAI21X1 OAI21X1_458 ( .A(new_wire_166), .B(_1604_), .C(_1632_), .Y(_1448_) );
INVX1 INVX1_205 ( .A(_1598_), .Y(_1605_) );
NAND2X1 NAND2X1_242 ( .A(AN), .B(new_wire_168), .Y(_1606_) );
OAI21X1 OAI21X1_459 ( .A(new_wire_168), .B(_1605_), .C(_1606_), .Y(_1450_) );
NAND2X1 NAND2X1_243 ( .A(HC), .B(new_wire_172), .Y(_1607_) );
OAI21X1 OAI21X1_460 ( .A(new_wire_172), .B(_1526_), .C(_1607_), .Y(_1449_) );
NAND2X1 NAND2X1_244 ( .A(new_wire_332), .B(new_wire_170), .Y(_1608_) );
AOI21X1 AOI21X1_131 ( .A(_1508_), .B(_1487_), .C(_1481_), .Y(_1609_) );
OAI21X1 OAI21X1_461 ( .A(_1476_), .B(_1507_), .C(_1508_), .Y(_1610_) );
OAI21X1 OAI21X1_462 ( .A(_1509_), .B(_1610_), .C(new_wire_12), .Y(_1611_) );
OAI21X1 OAI21X1_463 ( .A(_1609_), .B(_1611_), .C(_1608_), .Y(_1451__0_) );
NAND2X1 NAND2X1_245 ( .A(new_wire_346), .B(new_wire_172), .Y(_1612_) );
OAI21X1 OAI21X1_464 ( .A(new_wire_172), .B(_1517_), .C(_1612_), .Y(_1451__1_) );
NAND2X1 NAND2X1_246 ( .A(new_wire_359), .B(new_wire_170), .Y(_1613_) );
OAI21X1 OAI21X1_465 ( .A(new_wire_170), .B(_1523_), .C(_1613_), .Y(_1451__2_) );
NAND2X1 NAND2X1_247 ( .A(new_wire_353), .B(new_wire_170), .Y(_1614_) );
OAI21X1 OAI21X1_466 ( .A(new_wire_171), .B(_1587_), .C(_1614_), .Y(_1451__3_) );
NAND2X1 NAND2X1_248 ( .A(new_wire_314), .B(new_wire_171), .Y(_1615_) );
NOR2X1 NOR2X1_239 ( .A(_1593_), .B(_1592_), .Y(_1616_) );
OAI21X1 OAI21X1_467 ( .A(_1527_), .B(_1526_), .C(new_wire_12), .Y(_1617_) );
OAI21X1 OAI21X1_468 ( .A(_1616_), .B(_1617_), .C(_1615_), .Y(_1451__4_) );
NAND2X1 NAND2X1_249 ( .A(new_wire_297), .B(new_wire_173), .Y(_1618_) );
OAI21X1 OAI21X1_469 ( .A(new_wire_173), .B(_1600_), .C(_1618_), .Y(_1451__5_) );
NAND2X1 NAND2X1_250 ( .A(new_wire_327), .B(new_wire_166), .Y(_1619_) );
OAI21X1 OAI21X1_470 ( .A(new_wire_166), .B(_1602_), .C(_1619_), .Y(_1451__6_) );
NAND2X1 NAND2X1_251 ( .A(new_wire_322), .B(new_wire_167), .Y(_1620_) );
OAI21X1 OAI21X1_471 ( .A(new_wire_167), .B(_1605_), .C(_1620_), .Y(_1451__7_) );
AOI21X1 AOI21X1_132 ( .A(_1540_), .B(new_wire_609), .C(_1543_), .Y(_1621_) );
NAND2X1 NAND2X1_252 ( .A(ALU_BI7), .B(new_wire_168), .Y(_1622_) );
OAI21X1 OAI21X1_472 ( .A(new_wire_168), .B(_1621_), .C(_1622_), .Y(_1447_) );
NAND2X1 NAND2X1_253 ( .A(ALU_AI7), .B(new_wire_169), .Y(_1623_) );
OAI21X1 OAI21X1_473 ( .A(_1534_), .B(new_wire_169), .C(_1623_), .Y(_1446_) );
XOR2X1 XOR2X1_3 ( .A(ALU_BI7), .B(ALU_AI7), .Y(_1624_) );
XNOR2X1 XNOR2X1_9 ( .A(new_wire_336), .B(AN), .Y(_1625_) );
XNOR2X1 XNOR2X1_10 ( .A(_1624_), .B(_1625_), .Y(AV) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(new_wire_72), .D(_1448_), .Q(CO) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(new_wire_66), .D(_1450_), .Q(AN) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(new_wire_57), .D(_1449_), .Q(HC) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(new_wire_51), .D(_1451__0_), .Q(ADD_0_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(new_wire_60), .D(_1451__1_), .Q(ADD_1_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(new_wire_51), .D(_1451__2_), .Q(ADD_2_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(new_wire_60), .D(_1451__3_), .Q(ADD_3_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(new_wire_60), .D(_1451__4_), .Q(ADD_4_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(new_wire_57), .D(_1451__5_), .Q(ADD_5_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(new_wire_66), .D(_1451__6_), .Q(ADD_6_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(new_wire_72), .D(_1451__7_), .Q(ADD_7_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(new_wire_66), .D(_1447_), .Q(ALU_BI7) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(new_wire_66), .D(_1446_), .Q(ALU_AI7) );
BUFX2 new_buffer_1 ( .A(RDY_bF_buf8), .Y(new_wire_1) );
BUFX2 new_buffer_2 ( .A(RDY_bF_buf8), .Y(new_wire_2) );
BUFX2 new_buffer_3 ( .A(RDY_bF_buf8), .Y(new_wire_3) );
BUFX2 new_buffer_4 ( .A(RDY_bF_buf7), .Y(new_wire_4) );
BUFX2 new_buffer_5 ( .A(RDY_bF_buf7), .Y(new_wire_5) );
BUFX2 new_buffer_6 ( .A(RDY_bF_buf7), .Y(new_wire_6) );
BUFX2 new_buffer_7 ( .A(RDY_bF_buf6), .Y(new_wire_7) );
BUFX2 new_buffer_8 ( .A(RDY_bF_buf6), .Y(new_wire_8) );
BUFX2 new_buffer_9 ( .A(RDY_bF_buf6), .Y(new_wire_9) );
BUFX2 new_buffer_10 ( .A(RDY_bF_buf5), .Y(new_wire_10) );
BUFX2 new_buffer_11 ( .A(RDY_bF_buf5), .Y(new_wire_11) );
BUFX2 new_buffer_12 ( .A(RDY_bF_buf5), .Y(new_wire_12) );
BUFX2 new_buffer_13 ( .A(RDY_bF_buf4), .Y(new_wire_13) );
BUFX2 new_buffer_14 ( .A(RDY_bF_buf4), .Y(new_wire_14) );
BUFX2 new_buffer_15 ( .A(RDY_bF_buf4), .Y(new_wire_15) );
BUFX2 new_buffer_16 ( .A(RDY_bF_buf3), .Y(new_wire_16) );
BUFX2 new_buffer_17 ( .A(RDY_bF_buf3), .Y(new_wire_17) );
BUFX2 new_buffer_18 ( .A(RDY_bF_buf3), .Y(new_wire_18) );
BUFX2 new_buffer_19 ( .A(RDY_bF_buf2), .Y(new_wire_19) );
BUFX2 new_buffer_20 ( .A(RDY_bF_buf2), .Y(new_wire_20) );
BUFX2 new_buffer_21 ( .A(RDY_bF_buf2), .Y(new_wire_21) );
BUFX2 new_buffer_22 ( .A(RDY_bF_buf1), .Y(new_wire_22) );
BUFX2 new_buffer_23 ( .A(RDY_bF_buf1), .Y(new_wire_23) );
BUFX2 new_buffer_24 ( .A(RDY_bF_buf1), .Y(new_wire_24) );
BUFX2 new_buffer_25 ( .A(RDY_bF_buf0), .Y(new_wire_25) );
BUFX2 new_buffer_26 ( .A(RDY_bF_buf0), .Y(new_wire_26) );
BUFX2 new_buffer_27 ( .A(RDY_bF_buf0), .Y(new_wire_27) );
BUFX2 new_buffer_28 ( .A(_799_), .Y(new_wire_28) );
BUFX2 new_buffer_29 ( .A(_799_), .Y(new_wire_29) );
BUFX2 new_buffer_30 ( .A(_799__bF_buf4), .Y(new_wire_30) );
BUFX2 new_buffer_31 ( .A(_799__bF_buf4), .Y(new_wire_31) );
BUFX2 new_buffer_32 ( .A(_799__bF_buf3), .Y(new_wire_32) );
BUFX2 new_buffer_33 ( .A(_799__bF_buf3), .Y(new_wire_33) );
BUFX2 new_buffer_34 ( .A(_799__bF_buf2), .Y(new_wire_34) );
BUFX2 new_buffer_35 ( .A(_799__bF_buf2), .Y(new_wire_35) );
BUFX2 new_buffer_36 ( .A(_799__bF_buf1), .Y(new_wire_36) );
BUFX2 new_buffer_37 ( .A(_799__bF_buf1), .Y(new_wire_37) );
BUFX2 new_buffer_38 ( .A(_799__bF_buf0), .Y(new_wire_38) );
BUFX2 new_buffer_39 ( .A(_799__bF_buf0), .Y(new_wire_39) );
BUFX2 new_buffer_40 ( .A(clk_bF_buf11), .Y(new_wire_40) );
BUFX2 new_buffer_41 ( .A(clk_bF_buf11), .Y(new_wire_41) );
BUFX2 new_buffer_42 ( .A(clk_bF_buf11), .Y(new_wire_42) );
BUFX2 new_buffer_43 ( .A(clk_bF_buf10), .Y(new_wire_43) );
BUFX2 new_buffer_44 ( .A(clk_bF_buf10), .Y(new_wire_44) );
BUFX2 new_buffer_45 ( .A(clk_bF_buf10), .Y(new_wire_45) );
BUFX2 new_buffer_46 ( .A(clk_bF_buf9), .Y(new_wire_46) );
BUFX2 new_buffer_47 ( .A(clk_bF_buf9), .Y(new_wire_47) );
BUFX2 new_buffer_48 ( .A(clk_bF_buf9), .Y(new_wire_48) );
BUFX2 new_buffer_49 ( .A(clk_bF_buf8), .Y(new_wire_49) );
BUFX2 new_buffer_50 ( .A(clk_bF_buf8), .Y(new_wire_50) );
BUFX2 new_buffer_51 ( .A(clk_bF_buf8), .Y(new_wire_51) );
BUFX2 new_buffer_52 ( .A(clk_bF_buf7), .Y(new_wire_52) );
BUFX2 new_buffer_53 ( .A(clk_bF_buf7), .Y(new_wire_53) );
BUFX2 new_buffer_54 ( .A(clk_bF_buf7), .Y(new_wire_54) );
BUFX2 new_buffer_55 ( .A(clk_bF_buf6), .Y(new_wire_55) );
BUFX2 new_buffer_56 ( .A(clk_bF_buf6), .Y(new_wire_56) );
BUFX2 new_buffer_57 ( .A(clk_bF_buf6), .Y(new_wire_57) );
BUFX2 new_buffer_58 ( .A(clk_bF_buf5), .Y(new_wire_58) );
BUFX2 new_buffer_59 ( .A(clk_bF_buf5), .Y(new_wire_59) );
BUFX2 new_buffer_60 ( .A(clk_bF_buf5), .Y(new_wire_60) );
BUFX2 new_buffer_61 ( .A(clk_bF_buf4), .Y(new_wire_61) );
BUFX2 new_buffer_62 ( .A(clk_bF_buf4), .Y(new_wire_62) );
BUFX2 new_buffer_63 ( .A(clk_bF_buf4), .Y(new_wire_63) );
BUFX2 new_buffer_64 ( .A(clk_bF_buf3), .Y(new_wire_64) );
BUFX2 new_buffer_65 ( .A(clk_bF_buf3), .Y(new_wire_65) );
BUFX2 new_buffer_66 ( .A(clk_bF_buf3), .Y(new_wire_66) );
BUFX2 new_buffer_67 ( .A(clk_bF_buf2), .Y(new_wire_67) );
BUFX2 new_buffer_68 ( .A(clk_bF_buf2), .Y(new_wire_68) );
BUFX2 new_buffer_69 ( .A(clk_bF_buf2), .Y(new_wire_69) );
BUFX2 new_buffer_70 ( .A(clk_bF_buf1), .Y(new_wire_70) );
BUFX2 new_buffer_71 ( .A(clk_bF_buf1), .Y(new_wire_71) );
BUFX2 new_buffer_72 ( .A(clk_bF_buf1), .Y(new_wire_72) );
BUFX2 new_buffer_73 ( .A(clk_bF_buf0), .Y(new_wire_73) );
BUFX2 new_buffer_74 ( .A(clk_bF_buf0), .Y(new_wire_74) );
BUFX2 new_buffer_75 ( .A(clk_bF_buf0), .Y(new_wire_75) );
BUFX2 new_buffer_76 ( .A(_1101__bF_buf3), .Y(new_wire_76) );
BUFX2 new_buffer_77 ( .A(_1101__bF_buf3), .Y(new_wire_77) );
BUFX2 new_buffer_78 ( .A(_1101__bF_buf2), .Y(new_wire_78) );
BUFX2 new_buffer_79 ( .A(_1101__bF_buf2), .Y(new_wire_79) );
BUFX2 new_buffer_80 ( .A(_1101__bF_buf1), .Y(new_wire_80) );
BUFX2 new_buffer_81 ( .A(_1101__bF_buf1), .Y(new_wire_81) );
BUFX2 new_buffer_82 ( .A(_1101__bF_buf0), .Y(new_wire_82) );
BUFX2 new_buffer_83 ( .A(_1101__bF_buf0), .Y(new_wire_83) );
BUFX2 new_buffer_84 ( .A(_849_), .Y(new_wire_84) );
BUFX2 new_buffer_85 ( .A(_849_), .Y(new_wire_85) );
BUFX2 new_buffer_86 ( .A(_849__bF_buf4), .Y(new_wire_86) );
BUFX2 new_buffer_87 ( .A(_849__bF_buf4), .Y(new_wire_87) );
BUFX2 new_buffer_88 ( .A(_849__bF_buf3), .Y(new_wire_88) );
BUFX2 new_buffer_89 ( .A(_849__bF_buf3), .Y(new_wire_89) );
BUFX2 new_buffer_90 ( .A(_849__bF_buf2), .Y(new_wire_90) );
BUFX2 new_buffer_91 ( .A(_849__bF_buf2), .Y(new_wire_91) );
BUFX2 new_buffer_92 ( .A(_849__bF_buf1), .Y(new_wire_92) );
BUFX2 new_buffer_93 ( .A(_849__bF_buf1), .Y(new_wire_93) );
BUFX2 new_buffer_94 ( .A(_849__bF_buf0), .Y(new_wire_94) );
BUFX2 new_buffer_95 ( .A(_849__bF_buf0), .Y(new_wire_95) );
BUFX2 new_buffer_96 ( .A(_825_), .Y(new_wire_96) );
BUFX2 new_buffer_97 ( .A(_825_), .Y(new_wire_97) );
BUFX2 new_buffer_98 ( .A(_825__bF_buf4), .Y(new_wire_98) );
BUFX2 new_buffer_99 ( .A(_825__bF_buf4), .Y(new_wire_99) );
BUFX2 new_buffer_100 ( .A(_825__bF_buf3), .Y(new_wire_100) );
BUFX2 new_buffer_101 ( .A(_825__bF_buf3), .Y(new_wire_101) );
BUFX2 new_buffer_102 ( .A(_825__bF_buf2), .Y(new_wire_102) );
BUFX2 new_buffer_103 ( .A(_825__bF_buf2), .Y(new_wire_103) );
BUFX2 new_buffer_104 ( .A(_825__bF_buf1), .Y(new_wire_104) );
BUFX2 new_buffer_105 ( .A(_825__bF_buf1), .Y(new_wire_105) );
BUFX2 new_buffer_106 ( .A(_825__bF_buf0), .Y(new_wire_106) );
BUFX2 new_buffer_107 ( .A(_825__bF_buf0), .Y(new_wire_107) );
BUFX2 new_buffer_108 ( .A(_155__bF_buf3), .Y(new_wire_108) );
BUFX2 new_buffer_109 ( .A(_155__bF_buf3), .Y(new_wire_109) );
BUFX2 new_buffer_110 ( .A(_155__bF_buf2), .Y(new_wire_110) );
BUFX2 new_buffer_111 ( .A(_155__bF_buf2), .Y(new_wire_111) );
BUFX2 new_buffer_112 ( .A(_822_), .Y(new_wire_112) );
BUFX2 new_buffer_113 ( .A(_822_), .Y(new_wire_113) );
BUFX2 new_buffer_114 ( .A(_822__bF_buf4), .Y(new_wire_114) );
BUFX2 new_buffer_115 ( .A(_822__bF_buf4), .Y(new_wire_115) );
BUFX2 new_buffer_116 ( .A(_822__bF_buf3), .Y(new_wire_116) );
BUFX2 new_buffer_117 ( .A(_822__bF_buf3), .Y(new_wire_117) );
BUFX2 new_buffer_118 ( .A(_822__bF_buf2), .Y(new_wire_118) );
BUFX2 new_buffer_119 ( .A(_822__bF_buf2), .Y(new_wire_119) );
BUFX2 new_buffer_120 ( .A(_822__bF_buf1), .Y(new_wire_120) );
BUFX2 new_buffer_121 ( .A(_822__bF_buf1), .Y(new_wire_121) );
BUFX2 new_buffer_122 ( .A(_822__bF_buf0), .Y(new_wire_122) );
BUFX2 new_buffer_123 ( .A(_822__bF_buf0), .Y(new_wire_123) );
BUFX2 new_buffer_124 ( .A(_152__bF_buf3), .Y(new_wire_124) );
BUFX2 new_buffer_125 ( .A(_152__bF_buf3), .Y(new_wire_125) );
BUFX2 new_buffer_126 ( .A(_152__bF_buf2), .Y(new_wire_126) );
BUFX2 new_buffer_127 ( .A(_152__bF_buf2), .Y(new_wire_127) );
BUFX2 new_buffer_128 ( .A(_795_), .Y(new_wire_128) );
BUFX2 new_buffer_129 ( .A(_795_), .Y(new_wire_129) );
BUFX2 new_buffer_130 ( .A(_795__bF_buf4), .Y(new_wire_130) );
BUFX2 new_buffer_131 ( .A(_795__bF_buf4), .Y(new_wire_131) );
BUFX2 new_buffer_132 ( .A(_795__bF_buf3), .Y(new_wire_132) );
BUFX2 new_buffer_133 ( .A(_795__bF_buf3), .Y(new_wire_133) );
BUFX2 new_buffer_134 ( .A(_795__bF_buf2), .Y(new_wire_134) );
BUFX2 new_buffer_135 ( .A(_795__bF_buf2), .Y(new_wire_135) );
BUFX2 new_buffer_136 ( .A(_795__bF_buf1), .Y(new_wire_136) );
BUFX2 new_buffer_137 ( .A(_795__bF_buf1), .Y(new_wire_137) );
BUFX2 new_buffer_138 ( .A(_795__bF_buf0), .Y(new_wire_138) );
BUFX2 new_buffer_139 ( .A(_795__bF_buf0), .Y(new_wire_139) );
BUFX2 new_buffer_140 ( .A(_651_), .Y(new_wire_140) );
BUFX2 new_buffer_141 ( .A(_651_), .Y(new_wire_141) );
BUFX2 new_buffer_142 ( .A(_651__bF_buf4), .Y(new_wire_142) );
BUFX2 new_buffer_143 ( .A(_651__bF_buf4), .Y(new_wire_143) );
BUFX2 new_buffer_144 ( .A(_651__bF_buf3), .Y(new_wire_144) );
BUFX2 new_buffer_145 ( .A(_651__bF_buf3), .Y(new_wire_145) );
BUFX2 new_buffer_146 ( .A(_651__bF_buf2), .Y(new_wire_146) );
BUFX2 new_buffer_147 ( .A(_651__bF_buf2), .Y(new_wire_147) );
BUFX2 new_buffer_148 ( .A(_651__bF_buf1), .Y(new_wire_148) );
BUFX2 new_buffer_149 ( .A(_651__bF_buf1), .Y(new_wire_149) );
BUFX2 new_buffer_150 ( .A(_651__bF_buf0), .Y(new_wire_150) );
BUFX2 new_buffer_151 ( .A(_651__bF_buf0), .Y(new_wire_151) );
BUFX2 new_buffer_152 ( .A(_1070_), .Y(new_wire_152) );
BUFX2 new_buffer_153 ( .A(_1070_), .Y(new_wire_153) );
BUFX2 new_buffer_154 ( .A(_1070__bF_buf4), .Y(new_wire_154) );
BUFX2 new_buffer_155 ( .A(_1070__bF_buf4), .Y(new_wire_155) );
BUFX2 new_buffer_156 ( .A(_1070__bF_buf3), .Y(new_wire_156) );
BUFX2 new_buffer_157 ( .A(_1070__bF_buf3), .Y(new_wire_157) );
BUFX2 new_buffer_158 ( .A(_1070__bF_buf2), .Y(new_wire_158) );
BUFX2 new_buffer_159 ( .A(_1070__bF_buf2), .Y(new_wire_159) );
BUFX2 new_buffer_160 ( .A(_1070__bF_buf1), .Y(new_wire_160) );
BUFX2 new_buffer_161 ( .A(_1070__bF_buf1), .Y(new_wire_161) );
BUFX2 new_buffer_162 ( .A(_1070__bF_buf0), .Y(new_wire_162) );
BUFX2 new_buffer_163 ( .A(_1070__bF_buf0), .Y(new_wire_163) );
BUFX2 new_buffer_164 ( .A(_830__bF_buf3), .Y(new_wire_164) );
BUFX2 new_buffer_165 ( .A(_830__bF_buf3), .Y(new_wire_165) );
BUFX2 new_buffer_166 ( .A(_1631__bF_buf3), .Y(new_wire_166) );
BUFX2 new_buffer_167 ( .A(_1631__bF_buf3), .Y(new_wire_167) );
BUFX2 new_buffer_168 ( .A(_1631__bF_buf2), .Y(new_wire_168) );
BUFX2 new_buffer_169 ( .A(_1631__bF_buf2), .Y(new_wire_169) );
BUFX2 new_buffer_170 ( .A(_1631__bF_buf1), .Y(new_wire_170) );
BUFX2 new_buffer_171 ( .A(_1631__bF_buf1), .Y(new_wire_171) );
BUFX2 new_buffer_172 ( .A(_1631__bF_buf0), .Y(new_wire_172) );
BUFX2 new_buffer_173 ( .A(_1631__bF_buf0), .Y(new_wire_173) );
BUFX2 new_buffer_174 ( .A(_1017_), .Y(new_wire_174) );
BUFX2 new_buffer_175 ( .A(_1017_), .Y(new_wire_175) );
BUFX2 new_buffer_176 ( .A(_1017__bF_buf7), .Y(new_wire_176) );
BUFX2 new_buffer_177 ( .A(_1017__bF_buf7), .Y(new_wire_177) );
BUFX2 new_buffer_178 ( .A(_1017__bF_buf7), .Y(new_wire_178) );
BUFX2 new_buffer_179 ( .A(_1017__bF_buf6), .Y(new_wire_179) );
BUFX2 new_buffer_180 ( .A(_1017__bF_buf6), .Y(new_wire_180) );
BUFX2 new_buffer_181 ( .A(_1017__bF_buf6), .Y(new_wire_181) );
BUFX2 new_buffer_182 ( .A(_1017__bF_buf5), .Y(new_wire_182) );
BUFX2 new_buffer_183 ( .A(_1017__bF_buf5), .Y(new_wire_183) );
BUFX2 new_buffer_184 ( .A(_1017__bF_buf5), .Y(new_wire_184) );
BUFX2 new_buffer_185 ( .A(_1017__bF_buf4), .Y(new_wire_185) );
BUFX2 new_buffer_186 ( .A(_1017__bF_buf4), .Y(new_wire_186) );
BUFX2 new_buffer_187 ( .A(_1017__bF_buf3), .Y(new_wire_187) );
BUFX2 new_buffer_188 ( .A(_1017__bF_buf3), .Y(new_wire_188) );
BUFX2 new_buffer_189 ( .A(_1017__bF_buf2), .Y(new_wire_189) );
BUFX2 new_buffer_190 ( .A(_1017__bF_buf2), .Y(new_wire_190) );
BUFX2 new_buffer_191 ( .A(_1017__bF_buf1), .Y(new_wire_191) );
BUFX2 new_buffer_192 ( .A(_1017__bF_buf1), .Y(new_wire_192) );
BUFX2 new_buffer_193 ( .A(_1017__bF_buf0), .Y(new_wire_193) );
BUFX2 new_buffer_194 ( .A(_1017__bF_buf0), .Y(new_wire_194) );
BUFX2 new_buffer_195 ( .A(_859__bF_buf3), .Y(new_wire_195) );
BUFX2 new_buffer_196 ( .A(_859__bF_buf3), .Y(new_wire_196) );
BUFX2 new_buffer_197 ( .A(_859__bF_buf2), .Y(new_wire_197) );
BUFX2 new_buffer_198 ( .A(_859__bF_buf2), .Y(new_wire_198) );
BUFX2 new_buffer_199 ( .A(_859__bF_buf1), .Y(new_wire_199) );
BUFX2 new_buffer_200 ( .A(_859__bF_buf1), .Y(new_wire_200) );
BUFX2 new_buffer_201 ( .A(_148__bF_buf3), .Y(new_wire_201) );
BUFX2 new_buffer_202 ( .A(_148__bF_buf3), .Y(new_wire_202) );
BUFX2 new_buffer_203 ( .A(_815__bF_buf3), .Y(new_wire_203) );
BUFX2 new_buffer_204 ( .A(_815__bF_buf3), .Y(new_wire_204) );
BUFX2 new_buffer_205 ( .A(_815__bF_buf2), .Y(new_wire_205) );
BUFX2 new_buffer_206 ( .A(_815__bF_buf2), .Y(new_wire_206) );
BUFX2 new_buffer_207 ( .A(_815__bF_buf1), .Y(new_wire_207) );
BUFX2 new_buffer_208 ( .A(_815__bF_buf1), .Y(new_wire_208) );
BUFX2 new_buffer_209 ( .A(_815__bF_buf0), .Y(new_wire_209) );
BUFX2 new_buffer_210 ( .A(_815__bF_buf0), .Y(new_wire_210) );
BUFX2 new_buffer_211 ( .A(_812__bF_buf3), .Y(new_wire_211) );
BUFX2 new_buffer_212 ( .A(_812__bF_buf3), .Y(new_wire_212) );
BUFX2 new_buffer_213 ( .A(_812__bF_buf2), .Y(new_wire_213) );
BUFX2 new_buffer_214 ( .A(_812__bF_buf2), .Y(new_wire_214) );
BUFX2 new_buffer_215 ( .A(_812__bF_buf1), .Y(new_wire_215) );
BUFX2 new_buffer_216 ( .A(_812__bF_buf1), .Y(new_wire_216) );
BUFX2 new_buffer_217 ( .A(_812__bF_buf0), .Y(new_wire_217) );
BUFX2 new_buffer_218 ( .A(_812__bF_buf0), .Y(new_wire_218) );
BUFX2 new_buffer_219 ( .A(_809_), .Y(new_wire_219) );
BUFX2 new_buffer_220 ( .A(_809_), .Y(new_wire_220) );
BUFX2 new_buffer_221 ( .A(_809__bF_buf4), .Y(new_wire_221) );
BUFX2 new_buffer_222 ( .A(_809__bF_buf4), .Y(new_wire_222) );
BUFX2 new_buffer_223 ( .A(_809__bF_buf3), .Y(new_wire_223) );
BUFX2 new_buffer_224 ( .A(_809__bF_buf3), .Y(new_wire_224) );
BUFX2 new_buffer_225 ( .A(_809__bF_buf2), .Y(new_wire_225) );
BUFX2 new_buffer_226 ( .A(_809__bF_buf2), .Y(new_wire_226) );
BUFX2 new_buffer_227 ( .A(_809__bF_buf1), .Y(new_wire_227) );
BUFX2 new_buffer_228 ( .A(_809__bF_buf1), .Y(new_wire_228) );
BUFX2 new_buffer_229 ( .A(_809__bF_buf0), .Y(new_wire_229) );
BUFX2 new_buffer_230 ( .A(_809__bF_buf0), .Y(new_wire_230) );
BUFX2 new_buffer_231 ( .A(state_0_), .Y(new_wire_231) );
BUFX2 new_buffer_232 ( .A(state_0_), .Y(new_wire_232) );
BUFX2 new_buffer_233 ( .A(state_1_), .Y(new_wire_233) );
BUFX2 new_buffer_234 ( .A(state_1_), .Y(new_wire_234) );
BUFX2 new_buffer_235 ( .A(_789_), .Y(new_wire_235) );
BUFX2 new_buffer_236 ( .A(_789_), .Y(new_wire_236) );
BUFX2 new_buffer_237 ( .A(state_2_), .Y(new_wire_237) );
BUFX2 new_buffer_238 ( .A(state_2_), .Y(new_wire_238) );
BUFX2 new_buffer_239 ( .A(state_3_), .Y(new_wire_239) );
BUFX2 new_buffer_240 ( .A(state_3_), .Y(new_wire_240) );
BUFX2 new_buffer_241 ( .A(_792_), .Y(new_wire_241) );
BUFX2 new_buffer_242 ( .A(_792_), .Y(new_wire_242) );
BUFX2 new_buffer_243 ( .A(state_5_), .Y(new_wire_243) );
BUFX2 new_buffer_244 ( .A(state_5_), .Y(new_wire_244) );
BUFX2 new_buffer_245 ( .A(_794_), .Y(new_wire_245) );
BUFX2 new_buffer_246 ( .A(_794_), .Y(new_wire_246) );
BUFX2 new_buffer_247 ( .A(_794_), .Y(new_wire_247) );
BUFX2 new_buffer_248 ( .A(_794_), .Y(new_wire_248) );
BUFX2 new_buffer_249 ( .A(_796_), .Y(new_wire_249) );
BUFX2 new_buffer_250 ( .A(_796_), .Y(new_wire_250) );
BUFX2 new_buffer_251 ( .A(_798_), .Y(new_wire_251) );
BUFX2 new_buffer_252 ( .A(_798_), .Y(new_wire_252) );
BUFX2 new_buffer_253 ( .A(_798_), .Y(new_wire_253) );
BUFX2 new_buffer_254 ( .A(_798_), .Y(new_wire_254) );
BUFX2 new_buffer_255 ( .A(_802_), .Y(new_wire_255) );
BUFX2 new_buffer_256 ( .A(_802_), .Y(new_wire_256) );
BUFX2 new_buffer_257 ( .A(_805_), .Y(new_wire_257) );
BUFX2 new_buffer_258 ( .A(_805_), .Y(new_wire_258) );
BUFX2 new_buffer_259 ( .A(_807_), .Y(new_wire_259) );
BUFX2 new_buffer_260 ( .A(_807_), .Y(new_wire_260) );
BUFX2 new_buffer_261 ( .A(_808_), .Y(new_wire_261) );
BUFX2 new_buffer_262 ( .A(_808_), .Y(new_wire_262) );
BUFX2 new_buffer_263 ( .A(_808_), .Y(new_wire_263) );
BUFX2 new_buffer_264 ( .A(_808_), .Y(new_wire_264) );
BUFX2 new_buffer_265 ( .A(_810_), .Y(new_wire_265) );
BUFX2 new_buffer_266 ( .A(_810_), .Y(new_wire_266) );
BUFX2 new_buffer_267 ( .A(_814_), .Y(new_wire_267) );
BUFX2 new_buffer_268 ( .A(_814_), .Y(new_wire_268) );
BUFX2 new_buffer_269 ( .A(_817_), .Y(new_wire_269) );
BUFX2 new_buffer_270 ( .A(_817_), .Y(new_wire_270) );
BUFX2 new_buffer_271 ( .A(_817_), .Y(new_wire_271) );
BUFX2 new_buffer_272 ( .A(_819_), .Y(new_wire_272) );
BUFX2 new_buffer_273 ( .A(_819_), .Y(new_wire_273) );
BUFX2 new_buffer_274 ( .A(_819_), .Y(new_wire_274) );
BUFX2 new_buffer_275 ( .A(_819_), .Y(new_wire_275) );
BUFX2 new_buffer_276 ( .A(_820_), .Y(new_wire_276) );
BUFX2 new_buffer_277 ( .A(_820_), .Y(new_wire_277) );
BUFX2 new_buffer_278 ( .A(_820_), .Y(new_wire_278) );
BUFX2 new_buffer_279 ( .A(_824_), .Y(new_wire_279) );
BUFX2 new_buffer_280 ( .A(_824_), .Y(new_wire_280) );
BUFX2 new_buffer_281 ( .A(_824_), .Y(new_wire_281) );
BUFX2 new_buffer_282 ( .A(_824_), .Y(new_wire_282) );
BUFX2 new_buffer_283 ( .A(_833_), .Y(new_wire_283) );
BUFX2 new_buffer_284 ( .A(_833_), .Y(new_wire_284) );
BUFX2 new_buffer_285 ( .A(_834_), .Y(new_wire_285) );
BUFX2 new_buffer_286 ( .A(_834_), .Y(new_wire_286) );
BUFX2 new_buffer_287 ( .A(_838_), .Y(new_wire_287) );
BUFX2 new_buffer_288 ( .A(_838_), .Y(new_wire_288) );
BUFX2 new_buffer_289 ( .A(_843_), .Y(new_wire_289) );
BUFX2 new_buffer_290 ( .A(_843_), .Y(new_wire_290) );
BUFX2 new_buffer_291 ( .A(_843_), .Y(new_wire_291) );
BUFX2 new_buffer_292 ( .A(_843_), .Y(new_wire_292) );
BUFX2 new_buffer_293 ( .A(DIMUX_5_), .Y(new_wire_293) );
BUFX2 new_buffer_294 ( .A(DIMUX_5_), .Y(new_wire_294) );
BUFX2 new_buffer_295 ( .A(ADD_5_), .Y(new_wire_295) );
BUFX2 new_buffer_296 ( .A(ADD_5_), .Y(new_wire_296) );
BUFX2 new_buffer_297 ( .A(ADD_5_), .Y(new_wire_297) );
BUFX2 new_buffer_298 ( .A(_846_), .Y(new_wire_298) );
BUFX2 new_buffer_299 ( .A(_846_), .Y(new_wire_299) );
BUFX2 new_buffer_300 ( .A(_847_), .Y(new_wire_300) );
BUFX2 new_buffer_301 ( .A(_847_), .Y(new_wire_301) );
BUFX2 new_buffer_302 ( .A(_850_), .Y(new_wire_302) );
BUFX2 new_buffer_303 ( .A(_850_), .Y(new_wire_303) );
BUFX2 new_buffer_304 ( .A(_850_), .Y(new_wire_304) );
BUFX2 new_buffer_305 ( .A(_856_), .Y(new_wire_305) );
BUFX2 new_buffer_306 ( .A(_856_), .Y(new_wire_306) );
BUFX2 new_buffer_307 ( .A(_860_), .Y(new_wire_307) );
BUFX2 new_buffer_308 ( .A(_860_), .Y(new_wire_308) );
BUFX2 new_buffer_309 ( .A(_863_), .Y(new_wire_309) );
BUFX2 new_buffer_310 ( .A(_863_), .Y(new_wire_310) );
BUFX2 new_buffer_311 ( .A(_863_), .Y(new_wire_311) );
BUFX2 new_buffer_312 ( .A(ADD_4_), .Y(new_wire_312) );
BUFX2 new_buffer_313 ( .A(ADD_4_), .Y(new_wire_313) );
BUFX2 new_buffer_314 ( .A(ADD_4_), .Y(new_wire_314) );
BUFX2 new_buffer_315 ( .A(_870_), .Y(new_wire_315) );
BUFX2 new_buffer_316 ( .A(_870_), .Y(new_wire_316) );
BUFX2 new_buffer_317 ( .A(_870_), .Y(new_wire_317) );
BUFX2 new_buffer_318 ( .A(_872_), .Y(new_wire_318) );
BUFX2 new_buffer_319 ( .A(_872_), .Y(new_wire_319) );
BUFX2 new_buffer_320 ( .A(ADD_7_), .Y(new_wire_320) );
BUFX2 new_buffer_321 ( .A(ADD_7_), .Y(new_wire_321) );
BUFX2 new_buffer_322 ( .A(ADD_7_), .Y(new_wire_322) );
BUFX2 new_buffer_323 ( .A(_883_), .Y(new_wire_323) );
BUFX2 new_buffer_324 ( .A(_883_), .Y(new_wire_324) );
BUFX2 new_buffer_325 ( .A(ADD_6_), .Y(new_wire_325) );
BUFX2 new_buffer_326 ( .A(ADD_6_), .Y(new_wire_326) );
BUFX2 new_buffer_327 ( .A(ADD_6_), .Y(new_wire_327) );
BUFX2 new_buffer_328 ( .A(_893_), .Y(new_wire_328) );
BUFX2 new_buffer_329 ( .A(_893_), .Y(new_wire_329) );
BUFX2 new_buffer_330 ( .A(ADD_0_), .Y(new_wire_330) );
BUFX2 new_buffer_331 ( .A(ADD_0_), .Y(new_wire_331) );
BUFX2 new_buffer_332 ( .A(ADD_0_), .Y(new_wire_332) );
BUFX2 new_buffer_333 ( .A(_905_), .Y(new_wire_333) );
BUFX2 new_buffer_334 ( .A(_905_), .Y(new_wire_334) );
BUFX2 new_buffer_335 ( .A(CO), .Y(new_wire_335) );
BUFX2 new_buffer_336 ( .A(CO), .Y(new_wire_336) );
BUFX2 new_buffer_337 ( .A(_914_), .Y(new_wire_337) );
BUFX2 new_buffer_338 ( .A(_914_), .Y(new_wire_338) );
BUFX2 new_buffer_339 ( .A(_915_), .Y(new_wire_339) );
BUFX2 new_buffer_340 ( .A(_915_), .Y(new_wire_340) );
BUFX2 new_buffer_341 ( .A(_916_), .Y(new_wire_341) );
BUFX2 new_buffer_342 ( .A(_916_), .Y(new_wire_342) );
BUFX2 new_buffer_343 ( .A(_920_), .Y(new_wire_343) );
BUFX2 new_buffer_344 ( .A(_920_), .Y(new_wire_344) );
BUFX2 new_buffer_345 ( .A(ADD_1_), .Y(new_wire_345) );
BUFX2 new_buffer_346 ( .A(ADD_1_), .Y(new_wire_346) );
BUFX2 new_buffer_347 ( .A(_931_), .Y(new_wire_347) );
BUFX2 new_buffer_348 ( .A(_931_), .Y(new_wire_348) );
BUFX2 new_buffer_349 ( .A(_933_), .Y(new_wire_349) );
BUFX2 new_buffer_350 ( .A(_933_), .Y(new_wire_350) );
BUFX2 new_buffer_351 ( .A(ADD_3_), .Y(new_wire_351) );
BUFX2 new_buffer_352 ( .A(ADD_3_), .Y(new_wire_352) );
BUFX2 new_buffer_353 ( .A(ADD_3_), .Y(new_wire_353) );
BUFX2 new_buffer_354 ( .A(_944_), .Y(new_wire_354) );
BUFX2 new_buffer_355 ( .A(_944_), .Y(new_wire_355) );
BUFX2 new_buffer_356 ( .A(ADD_2_), .Y(new_wire_356) );
BUFX2 new_buffer_357 ( .A(ADD_2_), .Y(new_wire_357) );
BUFX2 new_buffer_358 ( .A(ADD_2_), .Y(new_wire_358) );
BUFX2 new_buffer_359 ( .A(ADD_2_), .Y(new_wire_359) );
BUFX2 new_buffer_360 ( .A(_956_), .Y(new_wire_360) );
BUFX2 new_buffer_361 ( .A(_956_), .Y(new_wire_361) );
BUFX2 new_buffer_362 ( .A(DIMUX_3_), .Y(new_wire_362) );
BUFX2 new_buffer_363 ( .A(DIMUX_3_), .Y(new_wire_363) );
BUFX2 new_buffer_364 ( .A(_972_), .Y(new_wire_364) );
BUFX2 new_buffer_365 ( .A(_972_), .Y(new_wire_365) );
BUFX2 new_buffer_366 ( .A(_978_), .Y(new_wire_366) );
BUFX2 new_buffer_367 ( .A(_978_), .Y(new_wire_367) );
BUFX2 new_buffer_368 ( .A(DIMUX_2_), .Y(new_wire_368) );
BUFX2 new_buffer_369 ( .A(DIMUX_2_), .Y(new_wire_369) );
BUFX2 new_buffer_370 ( .A(_983_), .Y(new_wire_370) );
BUFX2 new_buffer_371 ( .A(_983_), .Y(new_wire_371) );
BUFX2 new_buffer_372 ( .A(DIMUX_1_), .Y(new_wire_372) );
BUFX2 new_buffer_373 ( .A(DIMUX_1_), .Y(new_wire_373) );
BUFX2 new_buffer_374 ( .A(DIMUX_0_), .Y(new_wire_374) );
BUFX2 new_buffer_375 ( .A(DIMUX_0_), .Y(new_wire_375) );
BUFX2 new_buffer_376 ( .A(_1016_), .Y(new_wire_376) );
BUFX2 new_buffer_377 ( .A(_1016_), .Y(new_wire_377) );
BUFX2 new_buffer_378 ( .A(_1019_), .Y(new_wire_378) );
BUFX2 new_buffer_379 ( .A(_1019_), .Y(new_wire_379) );
BUFX2 new_buffer_380 ( .A(_1028_), .Y(new_wire_380) );
BUFX2 new_buffer_381 ( .A(_1028_), .Y(new_wire_381) );
BUFX2 new_buffer_382 ( .A(_1052_), .Y(new_wire_382) );
BUFX2 new_buffer_383 ( .A(_1052_), .Y(new_wire_383) );
BUFX2 new_buffer_384 ( .A(DIMUX_6_), .Y(new_wire_384) );
BUFX2 new_buffer_385 ( .A(DIMUX_6_), .Y(new_wire_385) );
BUFX2 new_buffer_386 ( .A(_1064_), .Y(new_wire_386) );
BUFX2 new_buffer_387 ( .A(_1064_), .Y(new_wire_387) );
BUFX2 new_buffer_388 ( .A(DIMUX_7_), .Y(new_wire_388) );
BUFX2 new_buffer_389 ( .A(DIMUX_7_), .Y(new_wire_389) );
BUFX2 new_buffer_390 ( .A(_1071_), .Y(new_wire_390) );
BUFX2 new_buffer_391 ( .A(_1071_), .Y(new_wire_391) );
BUFX2 new_buffer_392 ( .A(_1072_), .Y(new_wire_392) );
BUFX2 new_buffer_393 ( .A(_1072_), .Y(new_wire_393) );
BUFX2 new_buffer_394 ( .A(IRHOLD_valid), .Y(new_wire_394) );
BUFX2 new_buffer_395 ( .A(IRHOLD_valid), .Y(new_wire_395) );
BUFX2 new_buffer_396 ( .A(IRHOLD_valid), .Y(new_wire_396) );
BUFX2 new_buffer_397 ( .A(_1073_), .Y(new_wire_397) );
BUFX2 new_buffer_398 ( .A(_1073_), .Y(new_wire_398) );
BUFX2 new_buffer_399 ( .A(_1080_), .Y(new_wire_399) );
BUFX2 new_buffer_400 ( .A(_1080_), .Y(new_wire_400) );
BUFX2 new_buffer_401 ( .A(_1084_), .Y(new_wire_401) );
BUFX2 new_buffer_402 ( .A(_1084_), .Y(new_wire_402) );
BUFX2 new_buffer_403 ( .A(_1086_), .Y(new_wire_403) );
BUFX2 new_buffer_404 ( .A(_1086_), .Y(new_wire_404) );
BUFX2 new_buffer_405 ( .A(_1087_), .Y(new_wire_405) );
BUFX2 new_buffer_406 ( .A(_1087_), .Y(new_wire_406) );
BUFX2 new_buffer_407 ( .A(_1090_), .Y(new_wire_407) );
BUFX2 new_buffer_408 ( .A(_1090_), .Y(new_wire_408) );
BUFX2 new_buffer_409 ( .A(_1090_), .Y(new_wire_409) );
BUFX2 new_buffer_410 ( .A(_1090_), .Y(new_wire_410) );
BUFX2 new_buffer_411 ( .A(_1092_), .Y(new_wire_411) );
BUFX2 new_buffer_412 ( .A(_1092_), .Y(new_wire_412) );
BUFX2 new_buffer_413 ( .A(_1093_), .Y(new_wire_413) );
BUFX2 new_buffer_414 ( .A(_1093_), .Y(new_wire_414) );
BUFX2 new_buffer_415 ( .A(_1094_), .Y(new_wire_415) );
BUFX2 new_buffer_416 ( .A(_1094_), .Y(new_wire_416) );
BUFX2 new_buffer_417 ( .A(_1094_), .Y(new_wire_417) );
BUFX2 new_buffer_418 ( .A(_1100_), .Y(new_wire_418) );
BUFX2 new_buffer_419 ( .A(_1100_), .Y(new_wire_419) );
BUFX2 new_buffer_420 ( .A(_1100_), .Y(new_wire_420) );
BUFX2 new_buffer_421 ( .A(_1102_), .Y(new_wire_421) );
BUFX2 new_buffer_422 ( .A(_1102_), .Y(new_wire_422) );
BUFX2 new_buffer_423 ( .A(_1102_), .Y(new_wire_423) );
BUFX2 new_buffer_424 ( .A(_1102_), .Y(new_wire_424) );
BUFX2 new_buffer_425 ( .A(_1119_), .Y(new_wire_425) );
BUFX2 new_buffer_426 ( .A(_1119_), .Y(new_wire_426) );
BUFX2 new_buffer_427 ( .A(_1138_), .Y(new_wire_427) );
BUFX2 new_buffer_428 ( .A(_1138_), .Y(new_wire_428) );
BUFX2 new_buffer_429 ( .A(_1140_), .Y(new_wire_429) );
BUFX2 new_buffer_430 ( .A(_1140_), .Y(new_wire_430) );
BUFX2 new_buffer_431 ( .A(_1145_), .Y(new_wire_431) );
BUFX2 new_buffer_432 ( .A(_1145_), .Y(new_wire_432) );
BUFX2 new_buffer_433 ( .A(_1145_), .Y(new_wire_433) );
BUFX2 new_buffer_434 ( .A(_1155_), .Y(new_wire_434) );
BUFX2 new_buffer_435 ( .A(_1155_), .Y(new_wire_435) );
BUFX2 new_buffer_436 ( .A(_1161_), .Y(new_wire_436) );
BUFX2 new_buffer_437 ( .A(_1161_), .Y(new_wire_437) );
BUFX2 new_buffer_438 ( .A(_1171_), .Y(new_wire_438) );
BUFX2 new_buffer_439 ( .A(_1171_), .Y(new_wire_439) );
BUFX2 new_buffer_440 ( .A(_1178_), .Y(new_wire_440) );
BUFX2 new_buffer_441 ( .A(_1178_), .Y(new_wire_441) );
BUFX2 new_buffer_442 ( .A(_1178_), .Y(new_wire_442) );
BUFX2 new_buffer_443 ( .A(_1182_), .Y(new_wire_443) );
BUFX2 new_buffer_444 ( .A(_1182_), .Y(new_wire_444) );
BUFX2 new_buffer_445 ( .A(_1183_), .Y(new_wire_445) );
BUFX2 new_buffer_446 ( .A(_1183_), .Y(new_wire_446) );
BUFX2 new_buffer_447 ( .A(_1192_), .Y(new_wire_447) );
BUFX2 new_buffer_448 ( .A(_1192_), .Y(new_wire_448) );
BUFX2 new_buffer_449 ( .A(_1196_), .Y(new_wire_449) );
BUFX2 new_buffer_450 ( .A(_1196_), .Y(new_wire_450) );
BUFX2 new_buffer_451 ( .A(_1205_), .Y(new_wire_451) );
BUFX2 new_buffer_452 ( .A(_1205_), .Y(new_wire_452) );
BUFX2 new_buffer_453 ( .A(_1226_), .Y(new_wire_453) );
BUFX2 new_buffer_454 ( .A(_1226_), .Y(new_wire_454) );
BUFX2 new_buffer_455 ( .A(_1236_), .Y(new_wire_455) );
BUFX2 new_buffer_456 ( .A(_1236_), .Y(new_wire_456) );
BUFX2 new_buffer_457 ( .A(_1251_), .Y(new_wire_457) );
BUFX2 new_buffer_458 ( .A(_1251_), .Y(new_wire_458) );
BUFX2 new_buffer_459 ( .A(_1265_), .Y(new_wire_459) );
BUFX2 new_buffer_460 ( .A(_1265_), .Y(new_wire_460) );
BUFX2 new_buffer_461 ( .A(_1266_), .Y(new_wire_461) );
BUFX2 new_buffer_462 ( .A(_1266_), .Y(new_wire_462) );
BUFX2 new_buffer_463 ( .A(_1267_), .Y(new_wire_463) );
BUFX2 new_buffer_464 ( .A(_1267_), .Y(new_wire_464) );
BUFX2 new_buffer_465 ( .A(_1274_), .Y(new_wire_465) );
BUFX2 new_buffer_466 ( .A(_1274_), .Y(new_wire_466) );
BUFX2 new_buffer_467 ( .A(_1275_), .Y(new_wire_467) );
BUFX2 new_buffer_468 ( .A(_1275_), .Y(new_wire_468) );
BUFX2 new_buffer_469 ( .A(_1279_), .Y(new_wire_469) );
BUFX2 new_buffer_470 ( .A(_1279_), .Y(new_wire_470) );
BUFX2 new_buffer_471 ( .A(_1287_), .Y(new_wire_471) );
BUFX2 new_buffer_472 ( .A(_1287_), .Y(new_wire_472) );
BUFX2 new_buffer_473 ( .A(_1291_), .Y(new_wire_473) );
BUFX2 new_buffer_474 ( .A(_1291_), .Y(new_wire_474) );
BUFX2 new_buffer_475 ( .A(_1291_), .Y(new_wire_475) );
BUFX2 new_buffer_476 ( .A(_1294_), .Y(new_wire_476) );
BUFX2 new_buffer_477 ( .A(_1294_), .Y(new_wire_477) );
BUFX2 new_buffer_478 ( .A(_1298_), .Y(new_wire_478) );
BUFX2 new_buffer_479 ( .A(_1298_), .Y(new_wire_479) );
BUFX2 new_buffer_480 ( .A(_1300_), .Y(new_wire_480) );
BUFX2 new_buffer_481 ( .A(_1300_), .Y(new_wire_481) );
BUFX2 new_buffer_482 ( .A(cond_code_1_), .Y(new_wire_482) );
BUFX2 new_buffer_483 ( .A(cond_code_1_), .Y(new_wire_483) );
BUFX2 new_buffer_484 ( .A(_1323_), .Y(new_wire_484) );
BUFX2 new_buffer_485 ( .A(_1323_), .Y(new_wire_485) );
BUFX2 new_buffer_486 ( .A(_1358_), .Y(new_wire_486) );
BUFX2 new_buffer_487 ( .A(_1358_), .Y(new_wire_487) );
BUFX2 new_buffer_488 ( .A(_1388_), .Y(new_wire_488) );
BUFX2 new_buffer_489 ( .A(_1388_), .Y(new_wire_489) );
BUFX2 new_buffer_490 ( .A(_1389_), .Y(new_wire_490) );
BUFX2 new_buffer_491 ( .A(_1389_), .Y(new_wire_491) );
BUFX2 new_buffer_492 ( .A(_43_), .Y(new_wire_492) );
BUFX2 new_buffer_493 ( .A(_43_), .Y(new_wire_493) );
BUFX2 new_buffer_494 ( .A(_81_), .Y(new_wire_494) );
BUFX2 new_buffer_495 ( .A(_81_), .Y(new_wire_495) );
BUFX2 new_buffer_496 ( .A(_86_), .Y(new_wire_496) );
BUFX2 new_buffer_497 ( .A(_86_), .Y(new_wire_497) );
BUFX2 new_buffer_498 ( .A(_106_), .Y(new_wire_498) );
BUFX2 new_buffer_499 ( .A(_106_), .Y(new_wire_499) );
BUFX2 new_buffer_500 ( .A(_114_), .Y(new_wire_500) );
BUFX2 new_buffer_501 ( .A(_114_), .Y(new_wire_501) );
BUFX2 new_buffer_502 ( .A(_117_), .Y(new_wire_502) );
BUFX2 new_buffer_503 ( .A(_117_), .Y(new_wire_503) );
BUFX2 new_buffer_504 ( .A(BI_0_), .Y(new_wire_504) );
BUFX2 new_buffer_505 ( .A(BI_0_), .Y(new_wire_505) );
BUFX2 new_buffer_506 ( .A(BI_1_), .Y(new_wire_506) );
BUFX2 new_buffer_507 ( .A(BI_1_), .Y(new_wire_507) );
BUFX2 new_buffer_508 ( .A(_125_), .Y(new_wire_508) );
BUFX2 new_buffer_509 ( .A(_125_), .Y(new_wire_509) );
BUFX2 new_buffer_510 ( .A(_132_), .Y(new_wire_510) );
BUFX2 new_buffer_511 ( .A(_132_), .Y(new_wire_511) );
BUFX2 new_buffer_512 ( .A(_145_), .Y(new_wire_512) );
BUFX2 new_buffer_513 ( .A(_145_), .Y(new_wire_513) );
BUFX2 new_buffer_514 ( .A(_145_), .Y(new_wire_514) );
BUFX2 new_buffer_515 ( .A(_146_), .Y(new_wire_515) );
BUFX2 new_buffer_516 ( .A(_146_), .Y(new_wire_516) );
BUFX2 new_buffer_517 ( .A(_146_), .Y(new_wire_517) );
BUFX2 new_buffer_518 ( .A(_172_), .Y(new_wire_518) );
BUFX2 new_buffer_519 ( .A(_172_), .Y(new_wire_519) );
BUFX2 new_buffer_520 ( .A(_173_), .Y(new_wire_520) );
BUFX2 new_buffer_521 ( .A(_173_), .Y(new_wire_521) );
BUFX2 new_buffer_522 ( .A(_269_), .Y(new_wire_522) );
BUFX2 new_buffer_523 ( .A(_269_), .Y(new_wire_523) );
BUFX2 new_buffer_524 ( .A(alu_op_0_), .Y(new_wire_524) );
BUFX2 new_buffer_525 ( .A(alu_op_0_), .Y(new_wire_525) );
BUFX2 new_buffer_526 ( .A(alu_op_0_), .Y(new_wire_526) );
BUFX2 new_buffer_527 ( .A(alu_op_2_), .Y(new_wire_527) );
BUFX2 new_buffer_528 ( .A(alu_op_2_), .Y(new_wire_528) );
BUFX2 new_buffer_529 ( .A(alu_op_2_), .Y(new_wire_529) );
BUFX2 new_buffer_530 ( .A(alu_op_2_), .Y(new_wire_530) );
BUFX2 new_buffer_531 ( .A(alu_op_3_), .Y(new_wire_531) );
BUFX2 new_buffer_532 ( .A(alu_op_3_), .Y(new_wire_532) );
BUFX2 new_buffer_533 ( .A(alu_op_3_), .Y(new_wire_533) );
BUFX2 new_buffer_534 ( .A(_280_), .Y(new_wire_534) );
BUFX2 new_buffer_535 ( .A(_280_), .Y(new_wire_535) );
BUFX2 new_buffer_536 ( .A(_280_), .Y(new_wire_536) );
BUFX2 new_buffer_537 ( .A(_283_), .Y(new_wire_537) );
BUFX2 new_buffer_538 ( .A(_283_), .Y(new_wire_538) );
BUFX2 new_buffer_539 ( .A(_287_), .Y(new_wire_539) );
BUFX2 new_buffer_540 ( .A(_287_), .Y(new_wire_540) );
BUFX2 new_buffer_541 ( .A(_293_), .Y(new_wire_541) );
BUFX2 new_buffer_542 ( .A(_293_), .Y(new_wire_542) );
BUFX2 new_buffer_543 ( .A(D), .Y(new_wire_543) );
BUFX2 new_buffer_544 ( .A(D), .Y(new_wire_544) );
BUFX2 new_buffer_545 ( .A(_1175_), .Y(new_wire_545) );
BUFX2 new_buffer_546 ( .A(_1175_), .Y(new_wire_546) );
BUFX2 new_buffer_547 ( .A(plp), .Y(new_wire_547) );
BUFX2 new_buffer_548 ( .A(plp), .Y(new_wire_548) );
BUFX2 new_buffer_549 ( .A(_324_), .Y(new_wire_549) );
BUFX2 new_buffer_550 ( .A(_324_), .Y(new_wire_550) );
BUFX2 new_buffer_551 ( .A(_330_), .Y(new_wire_551) );
BUFX2 new_buffer_552 ( .A(_330_), .Y(new_wire_552) );
BUFX2 new_buffer_553 ( .A(alu_shift_right), .Y(new_wire_553) );
BUFX2 new_buffer_554 ( .A(alu_shift_right), .Y(new_wire_554) );
BUFX2 new_buffer_555 ( .A(alu_shift_right), .Y(new_wire_555) );
BUFX2 new_buffer_556 ( .A(alu_shift_right), .Y(new_wire_556) );
BUFX2 new_buffer_557 ( .A(_343_), .Y(new_wire_557) );
BUFX2 new_buffer_558 ( .A(_343_), .Y(new_wire_558) );
BUFX2 new_buffer_559 ( .A(_415_), .Y(new_wire_559) );
BUFX2 new_buffer_560 ( .A(_415_), .Y(new_wire_560) );
BUFX2 new_buffer_561 ( .A(_471_), .Y(new_wire_561) );
BUFX2 new_buffer_562 ( .A(_471_), .Y(new_wire_562) );
BUFX2 new_buffer_563 ( .A(_471_), .Y(new_wire_563) );
BUFX2 new_buffer_564 ( .A(_471_), .Y(new_wire_564) );
BUFX2 new_buffer_565 ( .A(_524_), .Y(new_wire_565) );
BUFX2 new_buffer_566 ( .A(_524_), .Y(new_wire_566) );
BUFX2 new_buffer_567 ( .A(_525_), .Y(new_wire_567) );
BUFX2 new_buffer_568 ( .A(_525_), .Y(new_wire_568) );
BUFX2 new_buffer_569 ( .A(_525_), .Y(new_wire_569) );
BUFX2 new_buffer_570 ( .A(_543_), .Y(new_wire_570) );
BUFX2 new_buffer_571 ( .A(_543_), .Y(new_wire_571) );
BUFX2 new_buffer_572 ( .A(_550_), .Y(new_wire_572) );
BUFX2 new_buffer_573 ( .A(_550_), .Y(new_wire_573) );
BUFX2 new_buffer_574 ( .A(_550_), .Y(new_wire_574) );
BUFX2 new_buffer_575 ( .A(_550_), .Y(new_wire_575) );
BUFX2 new_buffer_576 ( .A(_589_), .Y(new_wire_576) );
BUFX2 new_buffer_577 ( .A(_589_), .Y(new_wire_577) );
BUFX2 new_buffer_578 ( .A(_591_), .Y(new_wire_578) );
BUFX2 new_buffer_579 ( .A(_591_), .Y(new_wire_579) );
BUFX2 new_buffer_580 ( .A(_591_), .Y(new_wire_580) );
BUFX2 new_buffer_581 ( .A(_600_), .Y(new_wire_581) );
BUFX2 new_buffer_582 ( .A(_600_), .Y(new_wire_582) );
BUFX2 new_buffer_583 ( .A(_604_), .Y(new_wire_583) );
BUFX2 new_buffer_584 ( .A(_604_), .Y(new_wire_584) );
BUFX2 new_buffer_585 ( .A(_604_), .Y(new_wire_585) );
BUFX2 new_buffer_586 ( .A(_605_), .Y(new_wire_586) );
BUFX2 new_buffer_587 ( .A(_605_), .Y(new_wire_587) );
BUFX2 new_buffer_588 ( .A(_609_), .Y(new_wire_588) );
BUFX2 new_buffer_589 ( .A(_609_), .Y(new_wire_589) );
BUFX2 new_buffer_590 ( .A(_609_), .Y(new_wire_590) );
BUFX2 new_buffer_591 ( .A(_613_), .Y(new_wire_591) );
BUFX2 new_buffer_592 ( .A(_613_), .Y(new_wire_592) );
BUFX2 new_buffer_593 ( .A(_613_), .Y(new_wire_593) );
BUFX2 new_buffer_594 ( .A(_613_), .Y(new_wire_594) );
BUFX2 new_buffer_595 ( .A(_616_), .Y(new_wire_595) );
BUFX2 new_buffer_596 ( .A(_616_), .Y(new_wire_596) );
BUFX2 new_buffer_597 ( .A(_702_), .Y(new_wire_597) );
BUFX2 new_buffer_598 ( .A(_702_), .Y(new_wire_598) );
BUFX2 new_buffer_599 ( .A(_703_), .Y(new_wire_599) );
BUFX2 new_buffer_600 ( .A(_703_), .Y(new_wire_600) );
BUFX2 new_buffer_601 ( .A(_743_), .Y(new_wire_601) );
BUFX2 new_buffer_602 ( .A(_743_), .Y(new_wire_602) );
BUFX2 new_buffer_603 ( .A(_755_), .Y(new_wire_603) );
BUFX2 new_buffer_604 ( .A(_755_), .Y(new_wire_604) );
BUFX2 new_buffer_605 ( .A(_1633_), .Y(new_wire_605) );
BUFX2 new_buffer_606 ( .A(_1633_), .Y(new_wire_606) );
BUFX2 new_buffer_607 ( .A(_1634_), .Y(new_wire_607) );
BUFX2 new_buffer_608 ( .A(_1634_), .Y(new_wire_608) );
BUFX2 new_buffer_609 ( .A(_1634_), .Y(new_wire_609) );
BUFX2 new_buffer_610 ( .A(_1639_), .Y(new_wire_610) );
BUFX2 new_buffer_611 ( .A(_1639_), .Y(new_wire_611) );
BUFX2 new_buffer_612 ( .A(_1648_), .Y(new_wire_612) );
BUFX2 new_buffer_613 ( .A(_1648_), .Y(new_wire_613) );
BUFX2 new_buffer_614 ( .A(_1652_), .Y(new_wire_614) );
BUFX2 new_buffer_615 ( .A(_1652_), .Y(new_wire_615) );
BUFX2 new_buffer_616 ( .A(_1654_), .Y(new_wire_616) );
BUFX2 new_buffer_617 ( .A(_1654_), .Y(new_wire_617) );
endmodule
module testcase1 (in, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12 , out13, out14, out15, out16, out17, out18, out19, out20);
input in;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
wire vdd = 1'b1;
wire gnd = 1'b0;
INVX1 INVX1_0 ( .A(in), .Y(w1) );
INVX1 INVX1_1 ( .A(new_wire_1), .Y(out1) );
INVX1 INVX1_2 ( .A(new_wire_4), .Y(out2) );
INVX1 INVX1_3 ( .A(new_wire_2), .Y(out3) );
INVX1 INVX1_4 ( .A(new_wire_6), .Y(out4) );
BUFX2 new_buffer_1 ( .A(w1), .Y(new_wire_1) );
BUFX2 new_buffer_2 ( .A(new_wire_3), .Y(new_wire_2) );
INVX1 INVX1_0_clone_[1] ( .A(in), .Y(new_wire_3) );
BUFX2 new_buffer_1_clone_[2] ( .A(new_wire_5), .Y(new_wire_4) );
INVX1 INVX1_0_clone_[3] ( .A(in), .Y(new_wire_5) );
BUFX2 new_buffer_2_clone_[4] ( .A(new_wire_7), .Y(new_wire_6) );
INVX1 INVX1_0_clone_[1]_clone_[5] ( .A(in), .Y(new_wire_7) );
endmodule
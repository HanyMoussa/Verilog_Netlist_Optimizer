module cpu (clk, reset, DI, IRQ, NMI, RDY, AB, DO, WE);
input clk;
input reset;
input IRQ;
input NMI;
input RDY;
output WE;
input [7:0] DI;
output [15:0] AB;
output [7:0] DO;
wire vdd = 1'b1;
wire gnd = 1'b0;
BUFX4 BUFX4_1 ( .A(RDY), .Y(RDY_bF_buf8) );
BUFX4 BUFX4_2 ( .A(RDY), .Y(RDY_bF_buf7) );
BUFX4 BUFX4_3 ( .A(RDY), .Y(RDY_bF_buf6) );
BUFX4 BUFX4_4 ( .A(RDY), .Y(RDY_bF_buf5) );
BUFX4 BUFX4_5 ( .A(RDY), .Y(RDY_bF_buf4) );
BUFX4 BUFX4_6 ( .A(RDY), .Y(RDY_bF_buf3) );
BUFX4 BUFX4_7 ( .A(RDY), .Y(RDY_bF_buf2) );
BUFX4 BUFX4_8 ( .A(RDY), .Y(RDY_bF_buf1) );
BUFX4 BUFX4_9 ( .A(RDY), .Y(RDY_bF_buf0) );
BUFX4 BUFX4_10 ( .A(_799_), .Y(_799__bF_buf4) );
BUFX4 BUFX4_11 ( .A(_799_), .Y(_799__bF_buf3) );
BUFX4 BUFX4_12 ( .A(_799_), .Y(_799__bF_buf2) );
BUFX4 BUFX4_13 ( .A(_799_), .Y(_799__bF_buf1) );
BUFX4 BUFX4_14 ( .A(_799_), .Y(_799__bF_buf0) );
BUFX4 BUFX4_15 ( .A(clk), .Y(clk_bF_buf11) );
BUFX4 BUFX4_16 ( .A(clk), .Y(clk_bF_buf10) );
BUFX4 BUFX4_17 ( .A(clk), .Y(clk_bF_buf9) );
BUFX4 BUFX4_18 ( .A(clk), .Y(clk_bF_buf8) );
BUFX4 BUFX4_19 ( .A(clk), .Y(clk_bF_buf7) );
BUFX4 BUFX4_20 ( .A(clk), .Y(clk_bF_buf6) );
BUFX4 BUFX4_21 ( .A(clk), .Y(clk_bF_buf5) );
BUFX4 BUFX4_22 ( .A(clk), .Y(clk_bF_buf4) );
BUFX4 BUFX4_23 ( .A(clk), .Y(clk_bF_buf3) );
BUFX4 BUFX4_24 ( .A(clk), .Y(clk_bF_buf2) );
BUFX4 BUFX4_25 ( .A(clk), .Y(clk_bF_buf1) );
BUFX4 BUFX4_26 ( .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_27 ( .A(_1101_), .Y(_1101__bF_buf3) );
BUFX4 BUFX4_28 ( .A(_1101_), .Y(_1101__bF_buf2) );
BUFX4 BUFX4_29 ( .A(_1101_), .Y(_1101__bF_buf1) );
BUFX4 BUFX4_30 ( .A(_1101_), .Y(_1101__bF_buf0) );
BUFX4 BUFX4_31 ( .A(_849_), .Y(_849__bF_buf4) );
BUFX4 BUFX4_32 ( .A(_849_), .Y(_849__bF_buf3) );
BUFX4 BUFX4_33 ( .A(_849_), .Y(_849__bF_buf2) );
BUFX4 BUFX4_34 ( .A(_849_), .Y(_849__bF_buf1) );
BUFX4 BUFX4_35 ( .A(_849_), .Y(_849__bF_buf0) );
BUFX4 BUFX4_36 ( .A(_825_), .Y(_825__bF_buf4) );
BUFX4 BUFX4_37 ( .A(_825_), .Y(_825__bF_buf3) );
BUFX4 BUFX4_38 ( .A(_825_), .Y(_825__bF_buf2) );
BUFX4 BUFX4_39 ( .A(_825_), .Y(_825__bF_buf1) );
BUFX4 BUFX4_40 ( .A(_825_), .Y(_825__bF_buf0) );
BUFX4 BUFX4_41 ( .A(_822_), .Y(_822__bF_buf4) );
BUFX4 BUFX4_42 ( .A(_822_), .Y(_822__bF_buf3) );
BUFX4 BUFX4_43 ( .A(_822_), .Y(_822__bF_buf2) );
BUFX4 BUFX4_44 ( .A(_822_), .Y(_822__bF_buf1) );
BUFX4 BUFX4_45 ( .A(_822_), .Y(_822__bF_buf0) );
BUFX4 BUFX4_46 ( .A(_152_), .Y(_152__bF_buf3) );
BUFX4 BUFX4_47 ( .A(_152_), .Y(_152__bF_buf2) );
BUFX4 BUFX4_48 ( .A(_795_), .Y(_795__bF_buf4) );
BUFX4 BUFX4_49 ( .A(_795_), .Y(_795__bF_buf3) );
BUFX4 BUFX4_50 ( .A(_795_), .Y(_795__bF_buf2) );
BUFX4 BUFX4_51 ( .A(_795_), .Y(_795__bF_buf1) );
BUFX4 BUFX4_52 ( .A(_795_), .Y(_795__bF_buf0) );
BUFX4 BUFX4_53 ( .A(_651_), .Y(_651__bF_buf4) );
BUFX4 BUFX4_54 ( .A(_651_), .Y(_651__bF_buf3) );
BUFX4 BUFX4_55 ( .A(_651_), .Y(_651__bF_buf2) );
BUFX4 BUFX4_56 ( .A(_651_), .Y(_651__bF_buf1) );
BUFX4 BUFX4_57 ( .A(_651_), .Y(_651__bF_buf0) );
BUFX4 BUFX4_58 ( .A(_1070_), .Y(_1070__bF_buf4) );
BUFX4 BUFX4_59 ( .A(_1070_), .Y(_1070__bF_buf3) );
BUFX4 BUFX4_60 ( .A(_1070_), .Y(_1070__bF_buf2) );
BUFX4 BUFX4_61 ( .A(_1070_), .Y(_1070__bF_buf1) );
BUFX4 BUFX4_62 ( .A(_1070_), .Y(_1070__bF_buf0) );
BUFX4 BUFX4_63 ( .A(_1631_), .Y(_1631__bF_buf3) );
BUFX4 BUFX4_64 ( .A(_1631_), .Y(_1631__bF_buf2) );
BUFX4 BUFX4_65 ( .A(_1631_), .Y(_1631__bF_buf1) );
BUFX4 BUFX4_66 ( .A(_1631_), .Y(_1631__bF_buf0) );
BUFX4 BUFX4_67 ( .A(_1017_), .Y(_1017__bF_buf7) );
BUFX4 BUFX4_68 ( .A(_1017_), .Y(_1017__bF_buf6) );
BUFX4 BUFX4_69 ( .A(_1017_), .Y(_1017__bF_buf5) );
BUFX4 BUFX4_70 ( .A(_1017_), .Y(_1017__bF_buf4) );
BUFX4 BUFX4_71 ( .A(_1017_), .Y(_1017__bF_buf3) );
BUFX4 BUFX4_72 ( .A(_1017_), .Y(_1017__bF_buf2) );
BUFX4 BUFX4_73 ( .A(_1017_), .Y(_1017__bF_buf1) );
BUFX4 BUFX4_74 ( .A(_1017_), .Y(_1017__bF_buf0) );
BUFX4 BUFX4_75 ( .A(_859_), .Y(_859__bF_buf3) );
BUFX4 BUFX4_76 ( .A(_859_), .Y(_859__bF_buf2) );
BUFX4 BUFX4_77 ( .A(_148_), .Y(_148__bF_buf3) );
BUFX4 BUFX4_78 ( .A(_815_), .Y(_815__bF_buf3) );
BUFX4 BUFX4_79 ( .A(_815_), .Y(_815__bF_buf2) );
BUFX4 BUFX4_80 ( .A(_815_), .Y(_815__bF_buf1) );
BUFX4 BUFX4_81 ( .A(_815_), .Y(_815__bF_buf0) );
BUFX4 BUFX4_82 ( .A(_812_), .Y(_812__bF_buf3) );
BUFX4 BUFX4_83 ( .A(_812_), .Y(_812__bF_buf1) );
BUFX4 BUFX4_84 ( .A(_812_), .Y(_812__bF_buf0) );
BUFX4 BUFX4_85 ( .A(_809_), .Y(_809__bF_buf4) );
BUFX4 BUFX4_86 ( .A(_809_), .Y(_809__bF_buf3) );
BUFX4 BUFX4_87 ( .A(_809_), .Y(_809__bF_buf2) );
BUFX4 BUFX4_88 ( .A(_809_), .Y(_809__bF_buf1) );
BUFX4 BUFX4_89 ( .A(_809_), .Y(_809__bF_buf0) );
NAND2X1 NAND2X1_1 ( .A(state_0_), .B(state_1_), .Y(_788_) );
NOR2X1 NOR2X1_1 ( .A(state_3_), .B(_790_), .Y(_791_) );
NAND2X1 NAND2X1_2 ( .A(_789_), .B(_791_), .Y(_792_) );
NOR2X1 NOR2X1_2 ( .A(state_5_), .B(_793_), .Y(_794_) );
INVX8 INVX8_1 ( .A(_794_), .Y(_795_) );
NOR2X1 NOR2X1_3 ( .A(_795__bF_buf2), .B(_792_), .Y(_796_) );
NOR2X1 NOR2X1_4 ( .A(state_4_), .B(_797_), .Y(_798_) );
INVX8 INVX8_2 ( .A(_798_), .Y(_799_) );
NOR2X1 NOR2X1_5 ( .A(state_1_), .B(_800_), .Y(_801_) );
AND2X2 AND2X2_1 ( .A(state_2_), .B(state_3_), .Y(_802_) );
NAND2X1 NAND2X1_3 ( .A(_802_), .B(_801_), .Y(_803_) );
NOR2X1 NOR2X1_6 ( .A(state_2_), .B(_804_), .Y(_805_) );
NAND2X1 NAND2X1_4 ( .A(_801_), .B(_805_), .Y(_806_) );
AOI22X1 AOI22X1_1 ( .A(_795__bF_buf2), .B(_799__bF_buf1), .C(_803_), .D(_806_), .Y(_807_) );
NOR2X1 NOR2X1_7 ( .A(_796_), .B(_807_), .Y(_808_) );
OR2X2 OR2X2_1 ( .A(state_5_), .B(state_4_), .Y(_809_) );
NOR2X1 NOR2X1_8 ( .A(state_0_), .B(state_1_), .Y(_810_) );
NAND2X1 NAND2X1_5 ( .A(_810_), .B(_802_), .Y(_811_) );
NOR2X1 NOR2X1_9 ( .A(state_5_), .B(state_4_), .Y(_812_) );
NOR2X1 NOR2X1_10 ( .A(state_0_), .B(_813_), .Y(_814_) );
NAND3X1 NAND3X1_1 ( .A(_812__bF_buf0), .B(_791_), .C(_814_), .Y(_815_) );
OAI21X1 OAI21X1_1 ( .A(_809__bF_buf3), .B(_811_), .C(_815__bF_buf2), .Y(_816_) );
NAND3X1 NAND3X1_2 ( .A(_812__bF_buf1), .B(_805_), .C(_814_), .Y(_817_) );
OAI21X1 OAI21X1_2 ( .A(_809__bF_buf4), .B(_792_), .C(_817_), .Y(_818_) );
NOR2X1 NOR2X1_11 ( .A(_816_), .B(_818_), .Y(_819_) );
NAND2X1 NAND2X1_6 ( .A(_808_), .B(_819_), .Y(_820_) );
NAND3X1 NAND3X1_3 ( .A(_812__bF_buf0), .B(_810_), .C(_802_), .Y(_822_) );
INVX8 INVX8_3 ( .A(NMI_edge), .Y(_824_) );
OAI21X1 OAI21X1_3 ( .A(I), .B(_823_), .C(_824_), .Y(_825_) );
NOR2X1 NOR2X1_12 ( .A(_825__bF_buf4), .B(_822__bF_buf2), .Y(_826_) );
OAI21X1 OAI21X1_4 ( .A(_826_), .B(_821_), .C(PC_13_), .Y(_827_) );
NAND2X1 NAND2X1_7 ( .A(_823_), .B(_824_), .Y(_829_) );
OAI21X1 OAI21X1_5 ( .A(_828_), .B(NMI_edge), .C(_829_), .Y(_830_) );
NOR2X1 NOR2X1_13 ( .A(_822__bF_buf2), .B(_830__bF_buf0), .Y(_831_) );
NAND2X1 NAND2X1_8 ( .A(ABH_5_), .B(_831_), .Y(_832_) );
NAND2X1 NAND2X1_9 ( .A(state_2_), .B(_804_), .Y(_833_) );
NOR2X1 NOR2X1_14 ( .A(_788_), .B(_833_), .Y(_834_) );
NAND2X1 NAND2X1_10 ( .A(_794_), .B(_834_), .Y(_835_) );
NAND2X1 NAND2X1_11 ( .A(state_0_), .B(_813_), .Y(_836_) );
NAND2X1 NAND2X1_12 ( .A(state_2_), .B(state_3_), .Y(_837_) );
NOR2X1 NOR2X1_15 ( .A(_837_), .B(_836_), .Y(_838_) );
OAI21X1 OAI21X1_6 ( .A(_794_), .B(_798_), .C(_838_), .Y(_839_) );
NAND2X1 NAND2X1_13 ( .A(state_3_), .B(_790_), .Y(_840_) );
NOR2X1 NOR2X1_16 ( .A(_836_), .B(_840_), .Y(_841_) );
OAI21X1 OAI21X1_7 ( .A(_794_), .B(_798_), .C(_841_), .Y(_842_) );
NAND3X1 NAND3X1_4 ( .A(_835_), .B(_839_), .C(_842_), .Y(_843_) );
NAND2X1 NAND2X1_14 ( .A(RDY_bF_buf5), .B(DI[5]), .Y(_845_) );
OAI21X1 OAI21X1_8 ( .A(RDY_bF_buf5), .B(_844_), .C(_845_), .Y(DIMUX_5_) );
NAND3X1 NAND3X1_5 ( .A(_812__bF_buf1), .B(_789_), .C(_791_), .Y(_847_) );
NAND2X1 NAND2X1_15 ( .A(state_1_), .B(_800_), .Y(_848_) );
NOR3X1 NOR3X1_1 ( .A(_809__bF_buf4), .B(_833_), .C(_848_), .Y(_849_) );
NOR3X1 NOR3X1_2 ( .A(_809__bF_buf4), .B(_840_), .C(_848_), .Y(_850_) );
AOI21X1 AOI21X1_1 ( .A(_849__bF_buf2), .B(ABH_5_), .C(_850_), .Y(_851_) );
OAI21X1 OAI21X1_9 ( .A(_846_), .B(_847_), .C(_851_), .Y(_852_) );
AOI21X1 AOI21X1_2 ( .A(_843_), .B(DIMUX_5_), .C(_852_), .Y(_853_) );
NAND3X1 NAND3X1_6 ( .A(_832_), .B(_853_), .C(_827_), .Y(_854_) );
NAND3X1 NAND3X1_7 ( .A(PC_5_), .B(_808_), .C(_819_), .Y(_855_) );
NOR2X1 NOR2X1_17 ( .A(_840_), .B(_848_), .Y(_856_) );
AOI22X1 AOI22X1_2 ( .A(_812__bF_buf3), .B(_856_), .C(ADD_5_), .D(_849__bF_buf4), .Y(_857_) );
NAND3X1 NAND3X1_8 ( .A(PC_5_), .B(_812__bF_buf3), .C(_834_), .Y(_858_) );
INVX8 INVX8_4 ( .A(_822__bF_buf2), .Y(_859_) );
NOR2X1 NOR2X1_18 ( .A(_860_), .B(_825__bF_buf2), .Y(_861_) );
NAND2X1 NAND2X1_16 ( .A(IRQ), .B(_828_), .Y(_863_) );
AOI21X1 AOI21X1_3 ( .A(_863_), .B(_824_), .C(_862_), .Y(_864_) );
OAI21X1 OAI21X1_10 ( .A(_864_), .B(_861_), .C(_859__bF_buf3), .Y(_865_) );
NAND3X1 NAND3X1_9 ( .A(_858_), .B(_865_), .C(_857_), .Y(_866_) );
AOI21X1 AOI21X1_4 ( .A(ADD_5_), .B(_843_), .C(_866_), .Y(_867_) );
NAND3X1 NAND3X1_10 ( .A(PC_4_), .B(_808_), .C(_819_), .Y(_868_) );
AOI21X1 AOI21X1_5 ( .A(_849__bF_buf0), .B(ADD_4_), .C(_850_), .Y(_869_) );
NAND2X1 NAND2X1_17 ( .A(PC_4_), .B(_870_), .Y(_871_) );
NOR2X1 NOR2X1_19 ( .A(_872_), .B(_825__bF_buf2), .Y(_873_) );
AOI21X1 AOI21X1_6 ( .A(_863_), .B(_824_), .C(_874_), .Y(_875_) );
OAI21X1 OAI21X1_11 ( .A(_875_), .B(_873_), .C(_859__bF_buf3), .Y(_876_) );
NAND3X1 NAND3X1_11 ( .A(_876_), .B(_871_), .C(_869_), .Y(_877_) );
AOI21X1 AOI21X1_7 ( .A(ADD_4_), .B(_843_), .C(_877_), .Y(_878_) );
AOI22X1 AOI22X1_3 ( .A(_867_), .B(_855_), .C(_868_), .D(_878_), .Y(_879_) );
NAND3X1 NAND3X1_12 ( .A(PC_7_), .B(_808_), .C(_819_), .Y(_880_) );
AOI22X1 AOI22X1_4 ( .A(_812__bF_buf1), .B(_856_), .C(ADD_7_), .D(_849__bF_buf4), .Y(_881_) );
NAND3X1 NAND3X1_13 ( .A(PC_7_), .B(_812__bF_buf3), .C(_834_), .Y(_882_) );
NOR2X1 NOR2X1_20 ( .A(_883_), .B(_825__bF_buf4), .Y(_884_) );
AOI21X1 AOI21X1_8 ( .A(_863_), .B(_824_), .C(_885_), .Y(_886_) );
OAI21X1 OAI21X1_12 ( .A(_886_), .B(_884_), .C(_859__bF_buf0), .Y(_887_) );
NAND3X1 NAND3X1_14 ( .A(_882_), .B(_887_), .C(_881_), .Y(_888_) );
AOI21X1 AOI21X1_9 ( .A(ADD_7_), .B(_843_), .C(_888_), .Y(_889_) );
NAND3X1 NAND3X1_15 ( .A(PC_6_), .B(_808_), .C(_819_), .Y(_890_) );
AOI21X1 AOI21X1_10 ( .A(_849__bF_buf4), .B(ADD_6_), .C(_850_), .Y(_891_) );
NAND2X1 NAND2X1_18 ( .A(PC_6_), .B(_870_), .Y(_892_) );
NOR2X1 NOR2X1_21 ( .A(_893_), .B(_825__bF_buf4), .Y(_894_) );
AOI21X1 AOI21X1_11 ( .A(_863_), .B(_824_), .C(_895_), .Y(_896_) );
OAI21X1 OAI21X1_13 ( .A(_896_), .B(_894_), .C(_859__bF_buf0), .Y(_897_) );
NAND3X1 NAND3X1_16 ( .A(_897_), .B(_892_), .C(_891_), .Y(_898_) );
AOI21X1 AOI21X1_12 ( .A(ADD_6_), .B(_843_), .C(_898_), .Y(_899_) );
AOI22X1 AOI22X1_5 ( .A(_889_), .B(_880_), .C(_890_), .D(_899_), .Y(_900_) );
NAND2X1 NAND2X1_19 ( .A(_879_), .B(_900_), .Y(_901_) );
NAND3X1 NAND3X1_17 ( .A(PC_0_), .B(_808_), .C(_819_), .Y(_902_) );
OAI21X1 OAI21X1_14 ( .A(_796_), .B(_807_), .C(ADD_0_), .Y(_903_) );
OAI22X1 OAI22X1_1 ( .A(_905_), .B(_847_), .C(_904_), .D(_815__bF_buf0), .Y(_906_) );
NAND2X1 NAND2X1_20 ( .A(ABL_0_), .B(_825__bF_buf1), .Y(_907_) );
OAI21X1 OAI21X1_15 ( .A(_905_), .B(_825__bF_buf4), .C(_907_), .Y(_908_) );
AOI21X1 AOI21X1_13 ( .A(_859__bF_buf0), .B(_908_), .C(_906_), .Y(_909_) );
AND2X2 AND2X2_2 ( .A(_909_), .B(_903_), .Y(_910_) );
XOR2X1 XOR2X1_1 ( .A(CO), .B(backwards), .Y(_912_) );
OAI22X1 OAI22X1_2 ( .A(_822__bF_buf2), .B(_825__bF_buf4), .C(_912_), .D(_815__bF_buf1), .Y(_913_) );
NOR2X1 NOR2X1_22 ( .A(state_2_), .B(state_3_), .Y(_914_) );
NAND2X1 NAND2X1_21 ( .A(_914_), .B(_814_), .Y(_915_) );
NAND3X1 NAND3X1_18 ( .A(_789_), .B(_812__bF_buf1), .C(_805_), .Y(_916_) );
OAI21X1 OAI21X1_16 ( .A(_809__bF_buf4), .B(_915_), .C(_916_), .Y(_917_) );
NOR3X1 NOR3X1_3 ( .A(_917_), .B(_913_), .C(_911_), .Y(_918_) );
NAND2X1 NAND2X1_22 ( .A(_798_), .B(_838_), .Y(_919_) );
NOR2X1 NOR2X1_23 ( .A(_833_), .B(_836_), .Y(_920_) );
OAI21X1 OAI21X1_17 ( .A(_809__bF_buf4), .B(_921_), .C(_919_), .Y(_922_) );
NAND2X1 NAND2X1_23 ( .A(_810_), .B(_914_), .Y(_923_) );
OAI21X1 OAI21X1_18 ( .A(_838_), .B(_924_), .C(_812__bF_buf2), .Y(_925_) );
OAI21X1 OAI21X1_19 ( .A(state_5_), .B(_792_), .C(_925_), .Y(_926_) );
NOR2X1 NOR2X1_24 ( .A(_922_), .B(_926_), .Y(_927_) );
AOI22X1 AOI22X1_6 ( .A(_918_), .B(_927_), .C(_902_), .D(_910_), .Y(_928_) );
OAI21X1 OAI21X1_20 ( .A(_796_), .B(_807_), .C(ADD_1_), .Y(_929_) );
NAND3X1 NAND3X1_19 ( .A(PC_1_), .B(_808_), .C(_819_), .Y(_930_) );
OAI22X1 OAI22X1_3 ( .A(_931_), .B(_815__bF_buf0), .C(res), .D(_817_), .Y(_932_) );
NOR2X1 NOR2X1_25 ( .A(_933_), .B(_847_), .Y(_934_) );
NOR2X1 NOR2X1_26 ( .A(_934_), .B(_932_), .Y(_935_) );
NAND2X1 NAND2X1_24 ( .A(ABL_1_), .B(_825__bF_buf1), .Y(_936_) );
OAI21X1 OAI21X1_21 ( .A(_933_), .B(_825__bF_buf1), .C(_936_), .Y(_937_) );
NAND2X1 NAND2X1_25 ( .A(_859__bF_buf1), .B(_937_), .Y(_938_) );
AND2X2 AND2X2_3 ( .A(_935_), .B(_938_), .Y(_939_) );
NAND3X1 NAND3X1_20 ( .A(_929_), .B(_930_), .C(_939_), .Y(_940_) );
NAND3X1 NAND3X1_21 ( .A(PC_3_), .B(_808_), .C(_819_), .Y(_941_) );
AOI21X1 AOI21X1_14 ( .A(_849__bF_buf0), .B(ADD_3_), .C(_850_), .Y(_942_) );
NAND2X1 NAND2X1_26 ( .A(PC_3_), .B(_870_), .Y(_943_) );
NOR2X1 NOR2X1_27 ( .A(_944_), .B(_825__bF_buf2), .Y(_945_) );
AOI21X1 AOI21X1_15 ( .A(_863_), .B(_824_), .C(_946_), .Y(_947_) );
OAI21X1 OAI21X1_22 ( .A(_947_), .B(_945_), .C(_859__bF_buf3), .Y(_948_) );
NAND3X1 NAND3X1_22 ( .A(_948_), .B(_943_), .C(_942_), .Y(_949_) );
AOI21X1 AOI21X1_16 ( .A(ADD_3_), .B(_843_), .C(_949_), .Y(_950_) );
NAND3X1 NAND3X1_23 ( .A(PC_2_), .B(new_wire_33), .C(new_wire_35), .Y(_951_) );
NOR2X1 NOR2X1_28 ( .A(res), .B(_824_), .Y(_952_) );
AOI22X1 AOI22X1_7 ( .A(_849__bF_buf0), .B(ADD_2_), .C(_850_), .D(_953_), .Y(_954_) );
NAND2X1 NAND2X1_27 ( .A(PC_2_), .B(_870_), .Y(_955_) );
NOR2X1 NOR2X1_29 ( .A(_956_), .B(_825__bF_buf2), .Y(_957_) );
AOI21X1 AOI21X1_17 ( .A(_863_), .B(new_wire_40), .C(_958_), .Y(_959_) );
OAI21X1 OAI21X1_23 ( .A(_959_), .B(_957_), .C(_859__bF_buf3), .Y(_960_) );
NAND3X1 NAND3X1_24 ( .A(_955_), .B(_960_), .C(_954_), .Y(_961_) );
AOI21X1 AOI21X1_18 ( .A(ADD_2_), .B(_843_), .C(_961_), .Y(_962_) );
AOI22X1 AOI22X1_8 ( .A(_950_), .B(_941_), .C(_951_), .D(_962_), .Y(_963_) );
NAND3X1 NAND3X1_25 ( .A(_940_), .B(_928_), .C(_963_), .Y(_964_) );
NAND3X1 NAND3X1_26 ( .A(PC_11_), .B(new_wire_33), .C(new_wire_35), .Y(_965_) );
NAND2X1 NAND2X1_28 ( .A(RDY_bF_buf6), .B(DI[3]), .Y(_967_) );
OAI21X1 OAI21X1_24 ( .A(RDY_bF_buf6), .B(_966_), .C(_967_), .Y(DIMUX_3_) );
NAND3X1 NAND3X1_27 ( .A(ADD_3_), .B(_812__bF_buf3), .C(_834_), .Y(_968_) );
AOI21X1 AOI21X1_19 ( .A(_849__bF_buf3), .B(ABH_3_), .C(_850_), .Y(_969_) );
AOI21X1 AOI21X1_20 ( .A(_863_), .B(new_wire_40), .C(_970_), .Y(_971_) );
NOR2X1 NOR2X1_30 ( .A(_972_), .B(_825__bF_buf2), .Y(_973_) );
OAI21X1 OAI21X1_25 ( .A(_971_), .B(_973_), .C(_859__bF_buf1), .Y(_974_) );
NAND3X1 NAND3X1_28 ( .A(_968_), .B(_974_), .C(_969_), .Y(_975_) );
AOI21X1 AOI21X1_21 ( .A(_843_), .B(DIMUX_3_), .C(_975_), .Y(_976_) );
NAND3X1 NAND3X1_29 ( .A(PC_10_), .B(new_wire_33), .C(new_wire_35), .Y(_977_) );
MUX2X1 MUX2X1_1 ( .A(DI[2]), .B(DIHOLD_2_), .S(RDY_bF_buf5), .Y(_978_) );
NAND2X1 NAND2X1_29 ( .A(ADD_2_), .B(_870_), .Y(_979_) );
AOI21X1 AOI21X1_22 ( .A(_849__bF_buf1), .B(ABH_2_), .C(_850_), .Y(_980_) );
AOI21X1 AOI21X1_23 ( .A(_863_), .B(new_wire_40), .C(_981_), .Y(_982_) );
NOR2X1 NOR2X1_31 ( .A(_983_), .B(_825__bF_buf1), .Y(_984_) );
OAI21X1 OAI21X1_26 ( .A(_982_), .B(_984_), .C(_859__bF_buf1), .Y(_985_) );
NAND3X1 NAND3X1_30 ( .A(_985_), .B(_979_), .C(_980_), .Y(_986_) );
AOI21X1 AOI21X1_24 ( .A(new_wire_41), .B(DIMUX_2_), .C(_986_), .Y(_987_) );
AOI22X1 AOI22X1_9 ( .A(_976_), .B(_965_), .C(_977_), .D(_987_), .Y(_988_) );
NAND3X1 NAND3X1_31 ( .A(PC_9_), .B(new_wire_33), .C(new_wire_35), .Y(_989_) );
NAND2X1 NAND2X1_30 ( .A(RDY_bF_buf7), .B(DI[1]), .Y(_991_) );
OAI21X1 OAI21X1_27 ( .A(RDY_bF_buf7), .B(_990_), .C(_991_), .Y(DIMUX_1_) );
NAND3X1 NAND3X1_32 ( .A(ADD_1_), .B(_812__bF_buf3), .C(_834_), .Y(_992_) );
AOI21X1 AOI21X1_25 ( .A(_849__bF_buf0), .B(ABH_1_), .C(_850_), .Y(_993_) );
AOI21X1 AOI21X1_26 ( .A(new_wire_44), .B(new_wire_40), .C(_994_), .Y(_995_) );
NOR2X1 NOR2X1_32 ( .A(_996_), .B(_825__bF_buf2), .Y(_997_) );
OAI21X1 OAI21X1_28 ( .A(_995_), .B(_997_), .C(_859__bF_buf3), .Y(_998_) );
NAND3X1 NAND3X1_33 ( .A(_992_), .B(_998_), .C(_993_), .Y(_999_) );
AOI21X1 AOI21X1_27 ( .A(new_wire_41), .B(DIMUX_1_), .C(_999_), .Y(_1000_) );
NAND3X1 NAND3X1_34 ( .A(PC_8_), .B(new_wire_33), .C(new_wire_35), .Y(_1001_) );
NAND2X1 NAND2X1_31 ( .A(RDY_bF_buf5), .B(DI[0]), .Y(_1003_) );
OAI21X1 OAI21X1_29 ( .A(RDY_bF_buf5), .B(_1002_), .C(_1003_), .Y(DIMUX_0_) );
NAND2X1 NAND2X1_32 ( .A(ADD_0_), .B(_870_), .Y(_1004_) );
AOI21X1 AOI21X1_28 ( .A(_849__bF_buf0), .B(ABH_0_), .C(new_wire_43), .Y(_1005_) );
AOI21X1 AOI21X1_29 ( .A(new_wire_44), .B(new_wire_40), .C(_1006_), .Y(_1007_) );
NOR2X1 NOR2X1_33 ( .A(_1008_), .B(_825__bF_buf1), .Y(_1009_) );
OAI21X1 OAI21X1_30 ( .A(_1007_), .B(_1009_), .C(_859__bF_buf1), .Y(_1010_) );
NAND3X1 NAND3X1_35 ( .A(_1010_), .B(_1004_), .C(_1005_), .Y(_1011_) );
AOI21X1 AOI21X1_30 ( .A(new_wire_41), .B(DIMUX_0_), .C(_1011_), .Y(_1012_) );
AOI22X1 AOI22X1_10 ( .A(_1000_), .B(_989_), .C(_1001_), .D(_1012_), .Y(_1013_) );
NAND2X1 NAND2X1_33 ( .A(_988_), .B(_1013_), .Y(_1014_) );
NOR3X1 NOR3X1_4 ( .A(_901_), .B(_1014_), .C(_964_), .Y(_1015_) );
INVX8 INVX8_5 ( .A(RDY_bF_buf2), .Y(_1017_) );
OR2X2 OR2X2_2 ( .A(RDY_bF_buf5), .B(DIHOLD_4_), .Y(_1018_) );
OAI21X1 OAI21X1_31 ( .A(_1017__bF_buf4), .B(DI[4]), .C(_1018_), .Y(_1019_) );
OAI21X1 OAI21X1_32 ( .A(_1020_), .B(_815__bF_buf0), .C(_817_), .Y(_1021_) );
AOI21X1 AOI21X1_31 ( .A(ADD_4_), .B(_870_), .C(_1021_), .Y(_1022_) );
NOR2X1 NOR2X1_34 ( .A(_1016_), .B(_825__bF_buf1), .Y(_1023_) );
NOR2X1 NOR2X1_35 ( .A(_1020_), .B(_830__bF_buf0), .Y(_1024_) );
OAI21X1 OAI21X1_33 ( .A(_1023_), .B(_1024_), .C(_859__bF_buf1), .Y(_1025_) );
NAND2X1 NAND2X1_34 ( .A(_1025_), .B(_1022_), .Y(_1026_) );
AOI21X1 AOI21X1_32 ( .A(new_wire_41), .B(DIMUX_4_), .C(_1026_), .Y(_1027_) );
OAI21X1 OAI21X1_34 ( .A(_1016_), .B(_820_), .C(_1027_), .Y(_1028_) );
AOI21X1 AOI21X1_33 ( .A(_1015_), .B(_1028_), .C(_854_), .Y(_1029_) );
AND2X2 AND2X2_4 ( .A(_879_), .B(_900_), .Y(_1030_) );
NAND2X1 NAND2X1_35 ( .A(_940_), .B(_928_), .Y(_1031_) );
OAI21X1 OAI21X1_35 ( .A(_796_), .B(_807_), .C(ADD_3_), .Y(_1033_) );
AND2X2 AND2X2_5 ( .A(_942_), .B(_943_), .Y(_1034_) );
NAND3X1 NAND3X1_36 ( .A(_1033_), .B(_948_), .C(_1034_), .Y(_1035_) );
OAI21X1 OAI21X1_36 ( .A(_796_), .B(_807_), .C(ADD_2_), .Y(_1037_) );
AND2X2 AND2X2_6 ( .A(_954_), .B(_955_), .Y(_1038_) );
NAND3X1 NAND3X1_37 ( .A(_1037_), .B(_960_), .C(_1038_), .Y(_1039_) );
OAI22X1 OAI22X1_4 ( .A(_1035_), .B(_1032_), .C(_1036_), .D(_1039_), .Y(_1040_) );
NOR2X1 NOR2X1_36 ( .A(_1040_), .B(_1031_), .Y(_1041_) );
AND2X2 AND2X2_7 ( .A(_988_), .B(_1013_), .Y(_1042_) );
NAND3X1 NAND3X1_38 ( .A(_1030_), .B(_1042_), .C(_1041_), .Y(_1043_) );
NAND2X1 NAND2X1_36 ( .A(_1028_), .B(_854_), .Y(_1044_) );
OAI21X1 OAI21X1_37 ( .A(_1044_), .B(_1043_), .C(RDY_bF_buf3), .Y(_1045_) );
OAI22X1 OAI22X1_5 ( .A(_787_), .B(RDY_bF_buf5), .C(_1029_), .D(_1045_), .Y(_9__13_) );
NAND2X1 NAND2X1_37 ( .A(PC_14_), .B(_1017__bF_buf4), .Y(_1046_) );
NOR2X1 NOR2X1_37 ( .A(_1044_), .B(_1043_), .Y(_1047_) );
OAI21X1 OAI21X1_38 ( .A(_826_), .B(_821_), .C(PC_14_), .Y(_1048_) );
OAI21X1 OAI21X1_39 ( .A(_1049_), .B(_815__bF_buf0), .C(_817_), .Y(_1050_) );
AOI21X1 AOI21X1_34 ( .A(ADD_6_), .B(_870_), .C(_1050_), .Y(_1051_) );
MUX2X1 MUX2X1_2 ( .A(DI[6]), .B(DIHOLD_6_), .S(RDY_bF_buf0), .Y(_1052_) );
AOI22X1 AOI22X1_11 ( .A(ABH_6_), .B(_831_), .C(DIMUX_6_), .D(new_wire_41), .Y(_1053_) );
NAND3X1 NAND3X1_39 ( .A(_1051_), .B(_1053_), .C(_1048_), .Y(_1054_) );
NOR2X1 NOR2X1_38 ( .A(_1054_), .B(_1047_), .Y(_1055_) );
AND2X2 AND2X2_8 ( .A(_854_), .B(_1028_), .Y(_1056_) );
NAND3X1 NAND3X1_40 ( .A(_1056_), .B(_1054_), .C(_1015_), .Y(_1057_) );
NAND2X1 NAND2X1_38 ( .A(RDY_bF_buf3), .B(_1057_), .Y(_1058_) );
OAI21X1 OAI21X1_40 ( .A(_1058_), .B(_1055_), .C(_1046_), .Y(_9__14_) );
OAI21X1 OAI21X1_41 ( .A(_826_), .B(_821_), .C(PC_15_), .Y(_1060_) );
OAI21X1 OAI21X1_42 ( .A(_1061_), .B(_815__bF_buf0), .C(_817_), .Y(_1062_) );
AOI21X1 AOI21X1_35 ( .A(ABH_7_), .B(_831_), .C(_1062_), .Y(_1063_) );
MUX2X1 MUX2X1_3 ( .A(DI[7]), .B(DIHOLD_7_), .S(RDY_bF_buf5), .Y(_1064_) );
AOI22X1 AOI22X1_12 ( .A(ADD_7_), .B(new_wire_46), .C(DIMUX_7_), .D(new_wire_41), .Y(_1065_) );
NAND3X1 NAND3X1_41 ( .A(_1063_), .B(_1065_), .C(_1060_), .Y(_1066_) );
NAND3X1 NAND3X1_42 ( .A(_1054_), .B(_1067_), .C(_1047_), .Y(_1068_) );
AOI21X1 AOI21X1_36 ( .A(_1057_), .B(_1066_), .C(_1017__bF_buf4), .Y(_1069_) );
AOI22X1 AOI22X1_13 ( .A(_1017__bF_buf4), .B(_1059_), .C(_1068_), .D(_1069_), .Y(_9__15_) );
NOR2X1 NOR2X1_39 ( .A(_1017__bF_buf3), .B(_822__bF_buf0), .Y(_1070_) );
NAND2X1 NAND2X1_39 ( .A(_914_), .B(_801_), .Y(_1071_) );
NOR2X1 NOR2X1_40 ( .A(_799__bF_buf0), .B(_1071_), .Y(_1072_) );
NAND2X1 NAND2X1_40 ( .A(_1073_), .B(DIMUX_3_), .Y(_1075_) );
OAI21X1 OAI21X1_43 ( .A(_1073_), .B(_1074_), .C(_1075_), .Y(_1076_) );
NAND2X1 NAND2X1_41 ( .A(_830__bF_buf3), .B(_1076_), .Y(_1077_) );
NAND2X1 NAND2X1_42 ( .A(IRHOLD_valid), .B(IRHOLD_2_), .Y(_1078_) );
OAI21X1 OAI21X1_44 ( .A(IRHOLD_valid), .B(_978_), .C(_1078_), .Y(_1079_) );
AND2X2 AND2X2_9 ( .A(_1079_), .B(_830__bF_buf3), .Y(_1080_) );
NOR2X1 NOR2X1_41 ( .A(_1080_), .B(_1077_), .Y(_1081_) );
MUX2X1 MUX2X1_4 ( .A(DIMUX_1_), .B(IRHOLD_1_), .S(_1073_), .Y(_1082_) );
NOR2X1 NOR2X1_42 ( .A(_825__bF_buf3), .B(_1082_), .Y(_1083_) );
MUX2X1 MUX2X1_5 ( .A(DIMUX_0_), .B(IRHOLD_0_), .S(_1073_), .Y(_1084_) );
NOR2X1 NOR2X1_43 ( .A(_825__bF_buf3), .B(_1084_), .Y(_1085_) );
NOR2X1 NOR2X1_44 ( .A(_1083_), .B(_1085_), .Y(_1086_) );
NAND2X1 NAND2X1_43 ( .A(_1086_), .B(_1081_), .Y(_1087_) );
NAND2X1 NAND2X1_44 ( .A(IRHOLD_valid), .B(IRHOLD_7_), .Y(_1088_) );
OAI21X1 OAI21X1_45 ( .A(IRHOLD_valid), .B(_1064_), .C(_1088_), .Y(_1089_) );
NAND2X1 NAND2X1_45 ( .A(_830__bF_buf0), .B(_1089_), .Y(_1090_) );
NAND2X1 NAND2X1_46 ( .A(IRHOLD_valid), .B(IRHOLD_4_), .Y(_1091_) );
OAI21X1 OAI21X1_46 ( .A(IRHOLD_valid), .B(_1019_), .C(_1091_), .Y(_1092_) );
MUX2X1 MUX2X1_6 ( .A(DIMUX_5_), .B(IRHOLD_5_), .S(_1073_), .Y(_1093_) );
NOR2X1 NOR2X1_45 ( .A(_825__bF_buf0), .B(_1093_), .Y(_1094_) );
AOI21X1 AOI21X1_37 ( .A(_830__bF_buf2), .B(_1092_), .C(_1094_), .Y(_1095_) );
NAND2X1 NAND2X1_47 ( .A(_1090_), .B(_1095_), .Y(_1096_) );
NOR2X1 NOR2X1_46 ( .A(_1096_), .B(_1087_), .Y(_1097_) );
AOI22X1 AOI22X1_14 ( .A(_1017__bF_buf7), .B(_1072_), .C(_1070__bF_buf3), .D(_1097_), .Y(_1098_) );
NOR2X1 NOR2X1_47 ( .A(_809__bF_buf0), .B(_921_), .Y(_1099_) );
INVX8 INVX8_6 ( .A(_1070__bF_buf1), .Y(_1101_) );
AND2X2 AND2X2_10 ( .A(_1092_), .B(_830__bF_buf2), .Y(_1102_) );
OAI21X1 OAI21X1_47 ( .A(_1079_), .B(_1076_), .C(_830__bF_buf3), .Y(_1103_) );
NAND3X1 NAND3X1_43 ( .A(_1102_), .B(_1103_), .C(_1086_), .Y(_1104_) );
OAI22X1 OAI22X1_6 ( .A(RDY_bF_buf1), .B(_1100_), .C(_1101__bF_buf3), .D(_1104_), .Y(_1105_) );
NOR2X1 NOR2X1_48 ( .A(_836_), .B(_1106_), .Y(_1107_) );
NOR2X1 NOR2X1_49 ( .A(_797_), .B(_793_), .Y(_1108_) );
NAND2X1 NAND2X1_48 ( .A(_1108_), .B(_1107_), .Y(_1109_) );
NAND3X1 NAND3X1_44 ( .A(_810_), .B(_914_), .C(_1108_), .Y(_1110_) );
NAND2X1 NAND2X1_49 ( .A(RDY_bF_buf4), .B(_1111_), .Y(_1112_) );
OAI21X1 OAI21X1_48 ( .A(RDY_bF_buf4), .B(_1109_), .C(_1112_), .Y(_1113_) );
NAND2X1 NAND2X1_50 ( .A(_794_), .B(_1107_), .Y(_1114_) );
NAND2X1 NAND2X1_51 ( .A(_794_), .B(_924_), .Y(_1115_) );
MUX2X1 MUX2X1_7 ( .A(_1114_), .B(_1115_), .S(_1017__bF_buf0), .Y(_1116_) );
NOR2X1 NOR2X1_50 ( .A(_1116_), .B(_1113_), .Y(_1117_) );
OAI21X1 OAI21X1_49 ( .A(_799__bF_buf1), .B(_806_), .C(_1017__bF_buf0), .Y(_1118_) );
NAND2X1 NAND2X1_52 ( .A(_810_), .B(_805_), .Y(_1119_) );
OAI21X1 OAI21X1_50 ( .A(_799__bF_buf1), .B(_1119_), .C(RDY_bF_buf2), .Y(_1120_) );
AND2X2 AND2X2_11 ( .A(_1118_), .B(_1120_), .Y(_1121_) );
NAND2X1 NAND2X1_53 ( .A(_812__bF_buf2), .B(_841_), .Y(_1122_) );
NOR2X1 NOR2X1_51 ( .A(_809__bF_buf3), .B(_1119_), .Y(_1123_) );
NAND2X1 NAND2X1_54 ( .A(RDY_bF_buf8), .B(_1123_), .Y(_1124_) );
OAI21X1 OAI21X1_51 ( .A(RDY_bF_buf4), .B(_1122_), .C(_1124_), .Y(_1125_) );
NOR2X1 NOR2X1_52 ( .A(_1121_), .B(_1125_), .Y(_1126_) );
NOR2X1 NOR2X1_53 ( .A(_795__bF_buf2), .B(_1119_), .Y(_1127_) );
OAI21X1 OAI21X1_52 ( .A(_795__bF_buf2), .B(_806_), .C(_1017__bF_buf0), .Y(_1128_) );
OAI21X1 OAI21X1_53 ( .A(_1017__bF_buf0), .B(_1127_), .C(_1128_), .Y(_1129_) );
NOR2X1 NOR2X1_54 ( .A(_809__bF_buf0), .B(_1071_), .Y(_1130_) );
OAI21X1 OAI21X1_54 ( .A(_809__bF_buf0), .B(_923_), .C(RDY_bF_buf4), .Y(_1131_) );
OAI21X1 OAI21X1_55 ( .A(RDY_bF_buf4), .B(_1130_), .C(_1131_), .Y(_1132_) );
AND2X2 AND2X2_12 ( .A(_1129_), .B(_1132_), .Y(_1133_) );
NAND3X1 NAND3X1_45 ( .A(_1133_), .B(_1117_), .C(_1126_), .Y(_1134_) );
NOR2X1 NOR2X1_55 ( .A(_1134_), .B(_1105_), .Y(_1135_) );
OAI21X1 OAI21X1_56 ( .A(_1092_), .B(_1076_), .C(_830__bF_buf2), .Y(_1136_) );
NOR2X1 NOR2X1_56 ( .A(_788_), .B(_837_), .Y(_1137_) );
NOR2X1 NOR2X1_57 ( .A(_799__bF_buf2), .B(_1138_), .Y(_1139_) );
NAND2X1 NAND2X1_55 ( .A(_830__bF_buf3), .B(_1079_), .Y(_1140_) );
NOR2X1 NOR2X1_58 ( .A(_1140_), .B(_1101__bF_buf1), .Y(_1141_) );
AOI22X1 AOI22X1_15 ( .A(_1017__bF_buf7), .B(_1139_), .C(_1136_), .D(_1141_), .Y(_1142_) );
NAND2X1 NAND2X1_56 ( .A(_812__bF_buf2), .B(_1137_), .Y(_1143_) );
NAND2X1 NAND2X1_57 ( .A(_802_), .B(_814_), .Y(_1145_) );
OAI21X1 OAI21X1_57 ( .A(_809__bF_buf1), .B(_1145_), .C(RDY_bF_buf8), .Y(_1146_) );
OAI21X1 OAI21X1_58 ( .A(RDY_bF_buf8), .B(_1144_), .C(_1146_), .Y(_1147_) );
NAND2X1 NAND2X1_58 ( .A(_1147_), .B(_1142_), .Y(_1148_) );
NOR2X1 NOR2X1_59 ( .A(_833_), .B(_848_), .Y(_1149_) );
NAND2X1 NAND2X1_59 ( .A(_794_), .B(_1149_), .Y(_1150_) );
NAND2X1 NAND2X1_60 ( .A(RDY_bF_buf2), .B(_1150_), .Y(_1151_) );
OAI21X1 OAI21X1_59 ( .A(RDY_bF_buf2), .B(_796_), .C(_1151_), .Y(_1152_) );
NAND2X1 NAND2X1_61 ( .A(_798_), .B(_1149_), .Y(_1154_) );
NOR2X1 NOR2X1_60 ( .A(_799__bF_buf0), .B(_792_), .Y(_1155_) );
NAND2X1 NAND2X1_62 ( .A(_1017__bF_buf2), .B(_1155_), .Y(_1156_) );
OAI21X1 OAI21X1_60 ( .A(_1017__bF_buf2), .B(_1154_), .C(_1156_), .Y(_1157_) );
OR2X2 OR2X2_3 ( .A(_1153_), .B(_1157_), .Y(_1158_) );
NOR2X1 NOR2X1_61 ( .A(_1148_), .B(_1158_), .Y(_1159_) );
NAND2X1 NAND2X1_63 ( .A(_798_), .B(_856_), .Y(_1160_) );
NAND2X1 NAND2X1_64 ( .A(_789_), .B(_805_), .Y(_1161_) );
NOR2X1 NOR2X1_62 ( .A(_799__bF_buf1), .B(_1161_), .Y(_1162_) );
NAND2X1 NAND2X1_65 ( .A(_1017__bF_buf0), .B(_1162_), .Y(_1163_) );
OAI21X1 OAI21X1_61 ( .A(_1017__bF_buf0), .B(_1160_), .C(_1163_), .Y(_1164_) );
MUX2X1 MUX2X1_8 ( .A(_817_), .B(_916_), .S(RDY_bF_buf4), .Y(_1165_) );
OR2X2 OR2X2_4 ( .A(_1164_), .B(_1165_), .Y(_1166_) );
NAND2X1 NAND2X1_66 ( .A(RDY_bF_buf7), .B(_912_), .Y(_1167_) );
OAI22X1 OAI22X1_7 ( .A(RDY_bF_buf7), .B(_847_), .C(_815__bF_buf1), .D(_1167_), .Y(_1168_) );
NOR2X1 NOR2X1_63 ( .A(_795__bF_buf0), .B(_1161_), .Y(_1170_) );
NAND2X1 NAND2X1_67 ( .A(_805_), .B(_814_), .Y(_1171_) );
OAI21X1 OAI21X1_62 ( .A(_795__bF_buf0), .B(_1171_), .C(RDY_bF_buf2), .Y(_1172_) );
OAI21X1 OAI21X1_63 ( .A(RDY_bF_buf2), .B(_1170_), .C(_1172_), .Y(_1173_) );
NAND2X1 NAND2X1_68 ( .A(_1173_), .B(_1169_), .Y(_1174_) );
NOR2X1 NOR2X1_64 ( .A(_1174_), .B(_1166_), .Y(_1176_) );
NAND2X1 NAND2X1_69 ( .A(_1176_), .B(_1159_), .Y(_1177_) );
NAND2X1 NAND2X1_70 ( .A(_830__bF_buf1), .B(_1092_), .Y(_1178_) );
OAI21X1 OAI21X1_64 ( .A(_1073_), .B(IRHOLD_3_), .C(_830__bF_buf0), .Y(_1180_) );
AOI21X1 AOI21X1_38 ( .A(_1073_), .B(_1179_), .C(_1180_), .Y(_1181_) );
NAND2X1 NAND2X1_71 ( .A(_1140_), .B(_1181_), .Y(_1182_) );
OAI21X1 OAI21X1_65 ( .A(_825__bF_buf3), .B(_1082_), .C(_1085_), .Y(_1183_) );
NOR2X1 NOR2X1_65 ( .A(_1183_), .B(_1182_), .Y(_1184_) );
NAND2X1 NAND2X1_72 ( .A(_1178_), .B(_1184_), .Y(_1185_) );
NAND2X1 NAND2X1_73 ( .A(_1140_), .B(_1077_), .Y(_1186_) );
NOR2X1 NOR2X1_66 ( .A(_1090_), .B(_1102_), .Y(_1187_) );
OAI21X1 OAI21X1_66 ( .A(_825__bF_buf3), .B(_1084_), .C(_1187_), .Y(_1188_) );
OAI21X1 OAI21X1_67 ( .A(_1186_), .B(_1188_), .C(_1185_), .Y(_1189_) );
OAI21X1 OAI21X1_68 ( .A(_920_), .B(_1107_), .C(_794_), .Y(_1190_) );
NAND2X1 NAND2X1_74 ( .A(_798_), .B(_1191_), .Y(_1192_) );
NAND3X1 NAND3X1_46 ( .A(_839_), .B(_1190_), .C(_1192_), .Y(_1193_) );
OAI21X1 OAI21X1_69 ( .A(_809__bF_buf0), .B(_1071_), .C(_1109_), .Y(_1194_) );
NAND2X1 NAND2X1_75 ( .A(_800_), .B(_813_), .Y(_1195_) );
NOR2X1 NOR2X1_67 ( .A(_833_), .B(_1195_), .Y(_1196_) );
NAND2X1 NAND2X1_76 ( .A(_812__bF_buf0), .B(_1196_), .Y(_1197_) );
OAI21X1 OAI21X1_70 ( .A(_799__bF_buf0), .B(_1138_), .C(_1197_), .Y(_1198_) );
NOR2X1 NOR2X1_68 ( .A(_1198_), .B(_1194_), .Y(_1199_) );
NAND3X1 NAND3X1_47 ( .A(RDY_bF_buf8), .B(_1193_), .C(_1199_), .Y(_1200_) );
NAND3X1 NAND3X1_48 ( .A(_802_), .B(_810_), .C(_798_), .Y(_1201_) );
NAND2X1 NAND2X1_77 ( .A(RDY_bF_buf7), .B(_1202_), .Y(_1203_) );
OAI21X1 OAI21X1_71 ( .A(RDY_bF_buf7), .B(_919_), .C(_1203_), .Y(_1204_) );
NAND2X1 NAND2X1_78 ( .A(_812__bF_buf0), .B(_838_), .Y(_1205_) );
NAND2X1 NAND2X1_79 ( .A(new_wire_31), .B(_1196_), .Y(_1206_) );
NOR2X1 NOR2X1_69 ( .A(store), .B(CO), .Y(_1207_) );
NAND2X1 NAND2X1_80 ( .A(RDY_bF_buf0), .B(_1207_), .Y(_1208_) );
OAI22X1 OAI22X1_8 ( .A(RDY_bF_buf0), .B(_1205_), .C(_1208_), .D(_1206_), .Y(_1209_) );
NOR2X1 NOR2X1_70 ( .A(_788_), .B(_1106_), .Y(_1210_) );
NAND2X1 NAND2X1_81 ( .A(_812__bF_buf0), .B(_1210_), .Y(_1211_) );
AND2X2 AND2X2_13 ( .A(_1207_), .B(_1212_), .Y(_1213_) );
NAND2X1 NAND2X1_82 ( .A(RDY_bF_buf0), .B(_1213_), .Y(_1214_) );
NOR2X1 NOR2X1_71 ( .A(_1214_), .B(_1211_), .Y(_1215_) );
OR2X2 OR2X2_5 ( .A(_1215_), .B(_1209_), .Y(_1216_) );
NOR2X1 NOR2X1_72 ( .A(_1204_), .B(_1216_), .Y(_1217_) );
OR2X2 OR2X2_6 ( .A(_1194_), .B(_1198_), .Y(_1218_) );
NAND3X1 NAND3X1_49 ( .A(RDY_bF_buf1), .B(_1212_), .C(_1218_), .Y(_1219_) );
NAND3X1 NAND3X1_50 ( .A(_1200_), .B(_1219_), .C(_1217_), .Y(_1220_) );
AOI21X1 AOI21X1_39 ( .A(_1189_), .B(_1070__bF_buf4), .C(_1220_), .Y(_1221_) );
NAND2X1 NAND2X1_83 ( .A(_1103_), .B(_1086_), .Y(_1222_) );
OAI21X1 OAI21X1_72 ( .A(_1089_), .B(_1092_), .C(_830__bF_buf2), .Y(_1223_) );
NAND2X1 NAND2X1_84 ( .A(IRHOLD_valid), .B(IRHOLD_6_), .Y(_1224_) );
OAI21X1 OAI21X1_73 ( .A(new_wire_52), .B(_1052_), .C(_1224_), .Y(_1225_) );
NAND2X1 NAND2X1_85 ( .A(_830__bF_buf1), .B(_1225_), .Y(_1226_) );
NOR2X1 NOR2X1_73 ( .A(_1226_), .B(_1094_), .Y(_1227_) );
NAND2X1 NAND2X1_86 ( .A(_1223_), .B(_1227_), .Y(_1228_) );
NOR3X1 NOR3X1_5 ( .A(_1101__bF_buf1), .B(_1228_), .C(_1222_), .Y(_1229_) );
NAND3X1 NAND3X1_51 ( .A(_791_), .B(new_wire_32), .C(_801_), .Y(_1230_) );
NOR2X1 NOR2X1_74 ( .A(RDY_bF_buf4), .B(_1230_), .Y(_1231_) );
OAI21X1 OAI21X1_74 ( .A(_1207_), .B(_1206_), .C(RDY_bF_buf0), .Y(_1232_) );
OAI21X1 OAI21X1_75 ( .A(_795__bF_buf4), .B(_921_), .C(_1017__bF_buf2), .Y(_1233_) );
AND2X2 AND2X2_14 ( .A(_1232_), .B(_1233_), .Y(_1234_) );
NOR3X1 NOR3X1_6 ( .A(_1231_), .B(_1234_), .C(_1229_), .Y(_1235_) );
NAND2X1 NAND2X1_87 ( .A(_914_), .B(_789_), .Y(_1236_) );
NOR2X1 NOR2X1_75 ( .A(_1236_), .B(_799__bF_buf2), .Y(_1237_) );
NAND2X1 NAND2X1_88 ( .A(_1017__bF_buf6), .B(_1237_), .Y(_1238_) );
NAND3X1 NAND3X1_52 ( .A(RDY_bF_buf1), .B(write_back), .C(_1218_), .Y(_1239_) );
NOR2X1 NOR2X1_76 ( .A(_1236_), .B(_795__bF_buf1), .Y(_1240_) );
OAI21X1 OAI21X1_76 ( .A(_795__bF_buf1), .B(_915_), .C(RDY_bF_buf4), .Y(_1241_) );
OAI21X1 OAI21X1_77 ( .A(RDY_bF_buf8), .B(_1240_), .C(_1241_), .Y(_1242_) );
NAND3X1 NAND3X1_53 ( .A(_1238_), .B(_1242_), .C(_1239_), .Y(_1243_) );
NAND3X1 NAND3X1_54 ( .A(_802_), .B(_810_), .C(new_wire_31), .Y(_1244_) );
OAI21X1 OAI21X1_78 ( .A(_795__bF_buf0), .B(_803_), .C(_1017__bF_buf0), .Y(_1246_) );
OAI21X1 OAI21X1_79 ( .A(_1017__bF_buf0), .B(_1245_), .C(_1246_), .Y(_1247_) );
NOR2X1 NOR2X1_77 ( .A(_809__bF_buf1), .B(_915_), .Y(_1248_) );
OAI21X1 OAI21X1_80 ( .A(_809__bF_buf1), .B(_1236_), .C(_1017__bF_buf5), .Y(_1249_) );
OAI21X1 OAI21X1_81 ( .A(_1017__bF_buf5), .B(_1248_), .C(_1249_), .Y(_1250_) );
NOR2X1 NOR2X1_78 ( .A(_795__bF_buf4), .B(_1145_), .Y(_1251_) );
OAI21X1 OAI21X1_82 ( .A(_795__bF_buf1), .B(_1138_), .C(_1017__bF_buf5), .Y(_1252_) );
OAI21X1 OAI21X1_83 ( .A(_1017__bF_buf5), .B(_1251_), .C(_1252_), .Y(_1253_) );
NAND3X1 NAND3X1_55 ( .A(_1247_), .B(_1250_), .C(_1253_), .Y(_1254_) );
NOR2X1 NOR2X1_79 ( .A(_1254_), .B(_1243_), .Y(_1255_) );
NAND3X1 NAND3X1_56 ( .A(_1255_), .B(_1235_), .C(_1221_), .Y(_1256_) );
NOR2X1 NOR2X1_80 ( .A(_1177_), .B(_1256_), .Y(_1257_) );
NAND3X1 NAND3X1_57 ( .A(_1098_), .B(_1135_), .C(_1257_), .Y(_1438__0_) );
NAND3X1 NAND3X1_58 ( .A(_1250_), .B(_1253_), .C(_1258_), .Y(_1259_) );
NOR2X1 NOR2X1_81 ( .A(_1177_), .B(_1259_), .Y(_1260_) );
NAND2X1 NAND2X1_89 ( .A(_1017__bF_buf6), .B(_1251_), .Y(_1261_) );
AOI21X1 AOI21X1_40 ( .A(new_wire_52), .B(_1262_), .C(_825__bF_buf4), .Y(_1263_) );
OAI21X1 OAI21X1_84 ( .A(new_wire_52), .B(DIMUX_0_), .C(_1263_), .Y(_1264_) );
OAI21X1 OAI21X1_85 ( .A(_825__bF_buf4), .B(_1082_), .C(_1264_), .Y(_1265_) );
NOR2X1 NOR2X1_82 ( .A(_1265_), .B(_1182_), .Y(_1266_) );
AND2X2 AND2X2_15 ( .A(_1089_), .B(_830__bF_buf1), .Y(_1267_) );
NAND2X1 NAND2X1_90 ( .A(_1094_), .B(_1178_), .Y(_1268_) );
NOR2X1 NOR2X1_83 ( .A(_1267_), .B(_1268_), .Y(_1269_) );
NAND3X1 NAND3X1_59 ( .A(_1070__bF_buf1), .B(_1269_), .C(_1266_), .Y(_1270_) );
OAI21X1 OAI21X1_86 ( .A(_799__bF_buf2), .B(_1145_), .C(_1017__bF_buf6), .Y(_1271_) );
OAI21X1 OAI21X1_87 ( .A(_1017__bF_buf6), .B(_1237_), .C(_1271_), .Y(_1272_) );
NAND3X1 NAND3X1_60 ( .A(_1261_), .B(_1272_), .C(_1270_), .Y(_1273_) );
NAND2X1 NAND2X1_91 ( .A(_1090_), .B(_1178_), .Y(_1274_) );
AND2X2 AND2X2_16 ( .A(_1225_), .B(_830__bF_buf1), .Y(_1275_) );
OAI21X1 OAI21X1_88 ( .A(_825__bF_buf0), .B(_1093_), .C(_1275_), .Y(_1276_) );
NOR2X1 NOR2X1_84 ( .A(_1276_), .B(_1274_), .Y(_1277_) );
NAND2X1 NAND2X1_92 ( .A(_1080_), .B(_1181_), .Y(_1278_) );
NOR2X1 NOR2X1_85 ( .A(_1265_), .B(_1278_), .Y(_1279_) );
AND2X2 AND2X2_17 ( .A(_1279_), .B(_1277_), .Y(_1280_) );
OAI21X1 OAI21X1_89 ( .A(_795__bF_buf2), .B(_806_), .C(_916_), .Y(_1281_) );
NAND2X1 NAND2X1_93 ( .A(RDY_bF_buf2), .B(_1281_), .Y(_1282_) );
OAI21X1 OAI21X1_90 ( .A(RDY_bF_buf2), .B(_1150_), .C(_1282_), .Y(_1283_) );
AOI21X1 AOI21X1_41 ( .A(_1280_), .B(_1070__bF_buf4), .C(_1283_), .Y(_1284_) );
NOR2X1 NOR2X1_86 ( .A(_809__bF_buf1), .B(_1145_), .Y(_1285_) );
NAND2X1 NAND2X1_94 ( .A(_1017__bF_buf6), .B(_1285_), .Y(_1286_) );
NOR2X1 NOR2X1_87 ( .A(_1183_), .B(_1186_), .Y(_1287_) );
AND2X2 AND2X2_18 ( .A(_1287_), .B(_1178_), .Y(_1288_) );
NAND2X1 NAND2X1_95 ( .A(_1070__bF_buf4), .B(_1288_), .Y(_1289_) );
NAND3X1 NAND3X1_61 ( .A(_1286_), .B(_1289_), .C(_1284_), .Y(_1290_) );
NOR2X1 NOR2X1_88 ( .A(_795__bF_buf4), .B(_1171_), .Y(_1291_) );
NAND2X1 NAND2X1_96 ( .A(_1226_), .B(_1094_), .Y(_1292_) );
NAND2X1 NAND2X1_97 ( .A(_1223_), .B(_1293_), .Y(_1294_) );
NOR2X1 NOR2X1_89 ( .A(_1222_), .B(_1294_), .Y(_1295_) );
AOI22X1 AOI22X1_16 ( .A(_1017__bF_buf7), .B(_1291_), .C(_1070__bF_buf3), .D(_1295_), .Y(_1296_) );
NOR2X1 NOR2X1_90 ( .A(_1265_), .B(_1186_), .Y(_1298_) );
NAND2X1 NAND2X1_98 ( .A(_1275_), .B(_1094_), .Y(_1299_) );
NOR2X1 NOR2X1_91 ( .A(_1299_), .B(_1274_), .Y(_1300_) );
AND2X2 AND2X2_19 ( .A(_1298_), .B(_1300_), .Y(_1301_) );
AOI22X1 AOI22X1_17 ( .A(_1017__bF_buf7), .B(_1297_), .C(_1070__bF_buf3), .D(_1301_), .Y(_1302_) );
NAND2X1 NAND2X1_99 ( .A(cond_code_1_), .B(_1303_), .Y(_1304_) );
OAI21X1 OAI21X1_91 ( .A(cond_code_1_), .B(C), .C(_1304_), .Y(_1305_) );
NAND2X1 NAND2X1_100 ( .A(cond_code_1_), .B(_1306_), .Y(_1307_) );
OAI21X1 OAI21X1_92 ( .A(cond_code_1_), .B(N), .C(_1307_), .Y(_1308_) );
MUX2X1 MUX2X1_9 ( .A(_1305_), .B(_1308_), .S(cond_code_2_), .Y(_1309_) );
XNOR2X1 XNOR2X1_1 ( .A(_1309_), .B(cond_code_0_), .Y(_1310_) );
NAND3X1 NAND3X1_62 ( .A(RDY_bF_buf0), .B(_1099_), .C(_1310_), .Y(_1311_) );
NAND2X1 NAND2X1_101 ( .A(RDY_bF_buf7), .B(_1312_), .Y(_1313_) );
OAI21X1 OAI21X1_93 ( .A(new_wire_5), .B(_1154_), .C(_1313_), .Y(_1314_) );
AOI21X1 AOI21X1_42 ( .A(_1017__bF_buf2), .B(_849__bF_buf4), .C(_1314_), .Y(_1315_) );
AND2X2 AND2X2_20 ( .A(_1311_), .B(_1315_), .Y(_1316_) );
NAND3X1 NAND3X1_63 ( .A(_1316_), .B(_1302_), .C(_1296_), .Y(_1317_) );
NOR3X1 NOR3X1_7 ( .A(_1273_), .B(_1290_), .C(_1317_), .Y(_1318_) );
NAND2X1 NAND2X1_102 ( .A(new_wire_31), .B(_1319_), .Y(_1320_) );
OR2X2 OR2X2_7 ( .A(_1320_), .B(RDY_bF_buf1), .Y(_1321_) );
NAND3X1 NAND3X1_64 ( .A(_1102_), .B(_1070__bF_buf4), .C(_1287_), .Y(_1322_) );
NOR2X1 NOR2X1_92 ( .A(_799__bF_buf3), .B(_915_), .Y(_1323_) );
OAI21X1 OAI21X1_94 ( .A(_799__bF_buf0), .B(_1071_), .C(RDY_bF_buf8), .Y(_1324_) );
OAI21X1 OAI21X1_95 ( .A(RDY_bF_buf8), .B(_1323_), .C(_1324_), .Y(_1325_) );
NAND2X1 NAND2X1_103 ( .A(_1017__bF_buf2), .B(new_wire_43), .Y(_1326_) );
OAI21X1 OAI21X1_96 ( .A(_1017__bF_buf2), .B(_1122_), .C(_1326_), .Y(_1327_) );
AOI21X1 AOI21X1_43 ( .A(_1017__bF_buf5), .B(_1248_), .C(_1327_), .Y(_1328_) );
NAND2X1 NAND2X1_104 ( .A(_1325_), .B(_1328_), .Y(_1329_) );
OAI21X1 OAI21X1_97 ( .A(_1183_), .B(_1182_), .C(_1278_), .Y(_1330_) );
NOR2X1 NOR2X1_93 ( .A(_1101__bF_buf1), .B(_1178_), .Y(_1331_) );
AOI21X1 AOI21X1_44 ( .A(_1330_), .B(_1331_), .C(_1329_), .Y(_1332_) );
NAND3X1 NAND3X1_65 ( .A(_1321_), .B(_1322_), .C(_1332_), .Y(_1333_) );
NAND3X1 NAND3X1_66 ( .A(_1260_), .B(_1334_), .C(_1318_), .Y(_1438__1_) );
OAI21X1 OAI21X1_98 ( .A(_809__bF_buf1), .B(_811_), .C(_1017__bF_buf6), .Y(_1335_) );
NOR2X1 NOR2X1_94 ( .A(state_5_), .B(_792_), .Y(_1336_) );
AOI21X1 AOI21X1_45 ( .A(new_wire_32), .B(_841_), .C(_1336_), .Y(_1337_) );
NOR2X1 NOR2X1_95 ( .A(_1323_), .B(_1338_), .Y(_1339_) );
OAI21X1 OAI21X1_99 ( .A(_1196_), .B(_924_), .C(new_wire_32), .Y(_1340_) );
NAND3X1 NAND3X1_67 ( .A(_1340_), .B(_1337_), .C(_1339_), .Y(_1341_) );
NOR2X1 NOR2X1_96 ( .A(_912_), .B(_815__bF_buf1), .Y(_1342_) );
NOR2X1 NOR2X1_97 ( .A(_1017__bF_buf7), .B(_1342_), .Y(_1343_) );
OAI21X1 OAI21X1_100 ( .A(_1100_), .B(_1310_), .C(_1343_), .Y(_1344_) );
OR2X2 OR2X2_8 ( .A(_1344_), .B(_1341_), .Y(_1345_) );
NOR2X1 NOR2X1_98 ( .A(_1140_), .B(_1181_), .Y(_1346_) );
NOR2X1 NOR2X1_99 ( .A(_1101__bF_buf3), .B(_1346_), .Y(_1347_) );
OAI21X1 OAI21X1_101 ( .A(_1096_), .B(_1087_), .C(_1347_), .Y(_1348_) );
OAI21X1 OAI21X1_102 ( .A(_1102_), .B(_1277_), .C(_1298_), .Y(_1349_) );
NOR2X1 NOR2X1_100 ( .A(_1292_), .B(_1274_), .Y(_1350_) );
AOI22X1 AOI22X1_18 ( .A(_1279_), .B(_1277_), .C(_1298_), .D(_1350_), .Y(_1351_) );
AOI22X1 AOI22X1_19 ( .A(_1287_), .B(_1178_), .C(_1298_), .D(_1300_), .Y(_1352_) );
NAND3X1 NAND3X1_68 ( .A(_1349_), .B(_1351_), .C(_1352_), .Y(_1353_) );
NOR2X1 NOR2X1_101 ( .A(_1348_), .B(_1353_), .Y(_1354_) );
OAI21X1 OAI21X1_103 ( .A(_825__bF_buf3), .B(_1084_), .C(_1267_), .Y(_1355_) );
NOR2X1 NOR2X1_102 ( .A(_1102_), .B(_1355_), .Y(_1356_) );
AOI22X1 AOI22X1_20 ( .A(_1356_), .B(_1103_), .C(_1178_), .D(_1184_), .Y(_1357_) );
OAI21X1 OAI21X1_104 ( .A(_825__bF_buf3), .B(_1084_), .C(_1083_), .Y(_1358_) );
NOR2X1 NOR2X1_103 ( .A(_1358_), .B(_1182_), .Y(_1359_) );
AOI21X1 AOI21X1_46 ( .A(_1266_), .B(_1274_), .C(_1359_), .Y(_1360_) );
OR2X2 OR2X2_9 ( .A(_1093_), .B(_825__bF_buf0), .Y(_1361_) );
NOR2X1 NOR2X1_104 ( .A(_1267_), .B(_1361_), .Y(_1362_) );
NOR3X1 NOR3X1_8 ( .A(_1102_), .B(_1265_), .C(_1182_), .Y(_1363_) );
AOI22X1 AOI22X1_21 ( .A(_1102_), .B(_1330_), .C(_1362_), .D(_1363_), .Y(_1364_) );
NAND3X1 NAND3X1_69 ( .A(_1357_), .B(_1360_), .C(_1364_), .Y(_1365_) );
AOI21X1 AOI21X1_47 ( .A(_1292_), .B(_1090_), .C(_1102_), .Y(_1366_) );
NAND2X1 NAND2X1_105 ( .A(_1358_), .B(_1183_), .Y(_1367_) );
NOR2X1 NOR2X1_105 ( .A(new_wire_56), .B(_1278_), .Y(_1368_) );
AOI22X1 AOI22X1_22 ( .A(_1279_), .B(_1366_), .C(_1367_), .D(_1368_), .Y(_1369_) );
OAI21X1 OAI21X1_105 ( .A(_1089_), .B(_1225_), .C(_830__bF_buf3), .Y(_1370_) );
NAND3X1 NAND3X1_70 ( .A(_1095_), .B(_1370_), .C(_1298_), .Y(_1371_) );
AOI22X1 AOI22X1_23 ( .A(_1279_), .B(_1300_), .C(new_wire_56), .D(_1287_), .Y(_1372_) );
NAND3X1 NAND3X1_71 ( .A(_1371_), .B(_1369_), .C(_1372_), .Y(_1373_) );
NOR2X1 NOR2X1_106 ( .A(_1373_), .B(_1365_), .Y(_1374_) );
AOI22X1 AOI22X1_24 ( .A(_1335_), .B(_1345_), .C(_1354_), .D(_1374_), .Y(_1375_) );
OAI21X1 OAI21X1_106 ( .A(_795__bF_buf1), .B(_1376_), .C(_1017__bF_buf5), .Y(_1377_) );
OAI21X1 OAI21X1_107 ( .A(_1017__bF_buf5), .B(_1240_), .C(_1377_), .Y(_1378_) );
OAI21X1 OAI21X1_108 ( .A(_795__bF_buf0), .B(_1161_), .C(new_wire_5), .Y(_1380_) );
OAI21X1 OAI21X1_109 ( .A(new_wire_5), .B(_1245_), .C(_1380_), .Y(_1381_) );
OAI21X1 OAI21X1_110 ( .A(_799__bF_buf1), .B(_1161_), .C(new_wire_7), .Y(_1382_) );
OAI21X1 OAI21X1_111 ( .A(new_wire_7), .B(_1202_), .C(_1382_), .Y(_1383_) );
NAND2X1 NAND2X1_106 ( .A(_1383_), .B(_1381_), .Y(_1384_) );
NOR2X1 NOR2X1_107 ( .A(_1384_), .B(_1379_), .Y(_1385_) );
AND2X2 AND2X2_21 ( .A(_1375_), .B(_1385_), .Y(_1386_) );
OR2X2 OR2X2_10 ( .A(_1290_), .B(_1273_), .Y(_1387_) );
NAND2X1 NAND2X1_107 ( .A(_1081_), .B(_1388_), .Y(_1389_) );
OAI21X1 OAI21X1_112 ( .A(_1223_), .B(_1087_), .C(_1389_), .Y(_1390_) );
NAND2X1 NAND2X1_108 ( .A(_1070__bF_buf3), .B(_1390_), .Y(_1391_) );
NOR2X1 NOR2X1_108 ( .A(_799__bF_buf0), .B(_1376_), .Y(_1392_) );
NAND2X1 NAND2X1_109 ( .A(_1017__bF_buf6), .B(_1392_), .Y(_1393_) );
OAI21X1 OAI21X1_113 ( .A(_1213_), .B(_1211_), .C(RDY_bF_buf1), .Y(_1395_) );
OAI21X1 OAI21X1_114 ( .A(RDY_bF_buf1), .B(_1394_), .C(_1395_), .Y(_1396_) );
NAND3X1 NAND3X1_72 ( .A(_1393_), .B(_1396_), .C(_1391_), .Y(_1397_) );
NAND3X1 NAND3X1_73 ( .A(_1247_), .B(_1253_), .C(_1169_), .Y(_1398_) );
NOR2X1 NOR2X1_109 ( .A(_1398_), .B(_1105_), .Y(_1399_) );
NAND3X1 NAND3X1_74 ( .A(_1316_), .B(_1159_), .C(_1399_), .Y(_1400_) );
NOR2X1 NOR2X1_110 ( .A(_1397_), .B(_1400_), .Y(_1401_) );
NAND3X1 NAND3X1_75 ( .A(_1221_), .B(_1235_), .C(_1401_), .Y(_1402_) );
NOR2X1 NOR2X1_111 ( .A(_1387_), .B(_1402_), .Y(_1403_) );
NAND2X1 NAND2X1_110 ( .A(_1386_), .B(_1403_), .Y(_1438__2_) );
NAND3X1 NAND3X1_76 ( .A(_1070__bF_buf4), .B(_1300_), .C(_1279_), .Y(_1405_) );
OAI21X1 OAI21X1_115 ( .A(RDY_bF_buf1), .B(_1404_), .C(_1405_), .Y(_1406_) );
OAI21X1 OAI21X1_116 ( .A(_799__bF_buf2), .B(_1119_), .C(_1017__bF_buf5), .Y(_1407_) );
OAI21X1 OAI21X1_117 ( .A(_799__bF_buf2), .B(_792_), .C(RDY_bF_buf8), .Y(_1408_) );
AOI21X1 AOI21X1_48 ( .A(_1407_), .B(_1408_), .C(_1406_), .Y(_1409_) );
AOI22X1 AOI22X1_25 ( .A(_1017__bF_buf6), .B(_1111_), .C(_1331_), .D(_1346_), .Y(_1411_) );
OAI21X1 OAI21X1_118 ( .A(_923_), .B(_795__bF_buf1), .C(new_wire_28), .Y(_1412_) );
OAI21X1 OAI21X1_119 ( .A(new_wire_25), .B(_1144_), .C(_1412_), .Y(_1413_) );
NAND2X1 NAND2X1_111 ( .A(_1413_), .B(_1411_), .Y(_1414_) );
NAND2X1 NAND2X1_112 ( .A(_812__bF_buf2), .B(_924_), .Y(_1415_) );
NOR2X1 NOR2X1_112 ( .A(_923_), .B(_799__bF_buf2), .Y(_1416_) );
OAI21X1 OAI21X1_120 ( .A(_795__bF_buf4), .B(_1138_), .C(new_wire_1), .Y(_1417_) );
OAI21X1 OAI21X1_121 ( .A(new_wire_1), .B(_1416_), .C(_1417_), .Y(_1418_) );
OAI21X1 OAI21X1_122 ( .A(new_wire_1), .B(_1415_), .C(_1418_), .Y(_1419_) );
NOR2X1 NOR2X1_113 ( .A(_1419_), .B(_1414_), .Y(_1420_) );
OAI21X1 OAI21X1_123 ( .A(_1101__bF_buf3), .B(_1369_), .C(_1420_), .Y(_1421_) );
NOR2X1 NOR2X1_114 ( .A(_1421_), .B(_1410_), .Y(_1422_) );
NAND2X1 NAND2X1_113 ( .A(_1098_), .B(_1135_), .Y(_1423_) );
NOR3X1 NOR3X1_9 ( .A(_1333_), .B(_1397_), .C(_1423_), .Y(_1424_) );
NAND3X1 NAND3X1_77 ( .A(_1422_), .B(_1424_), .C(_1318_), .Y(_1425_) );
NAND3X1 NAND3X1_78 ( .A(_1385_), .B(_1375_), .C(_1257_), .Y(_1426_) );
OAI21X1 OAI21X1_124 ( .A(_1341_), .B(_1344_), .C(_1335_), .Y(_1427_) );
NAND2X1 NAND2X1_114 ( .A(_1354_), .B(_1374_), .Y(_1428_) );
NAND2X1 NAND2X1_115 ( .A(_1427_), .B(_1428_), .Y(_1429_) );
NAND2X1 NAND2X1_116 ( .A(_1178_), .B(_1287_), .Y(_1430_) );
OAI21X1 OAI21X1_125 ( .A(_1101__bF_buf3), .B(_1430_), .C(_1286_), .Y(_1431_) );
NAND2X1 NAND2X1_117 ( .A(_1173_), .B(_1253_), .Y(_1432_) );
NAND2X1 NAND2X1_118 ( .A(_1247_), .B(_1129_), .Y(_1433_) );
NOR2X1 NOR2X1_115 ( .A(_1433_), .B(_1432_), .Y(_1434_) );
OR2X2 OR2X2_11 ( .A(_1125_), .B(_1121_), .Y(_1435_) );
NOR2X1 NOR2X1_116 ( .A(_1327_), .B(_1435_), .Y(_1436_) );
NOR2X1 NOR2X1_117 ( .A(_1384_), .B(_1166_), .Y(_1437_) );
NAND3X1 NAND3X1_79 ( .A(_1434_), .B(_1437_), .C(_1436_), .Y(_41_) );
NOR3X1 NOR3X1_10 ( .A(_1148_), .B(_1431_), .C(_41_), .Y(_42_) );
NAND2X1 NAND2X1_119 ( .A(_1350_), .B(_1298_), .Y(_44_) );
OAI22X1 OAI22X1_9 ( .A(RDY_bF_buf1), .B(_43_), .C(_1101__bF_buf3), .D(_44_), .Y(_45_) );
NAND2X1 NAND2X1_120 ( .A(_1300_), .B(_1298_), .Y(_46_) );
OAI22X1 OAI22X1_10 ( .A(new_wire_8), .B(_1160_), .C(_1101__bF_buf3), .D(_46_), .Y(_47_) );
NOR3X1 NOR3X1_11 ( .A(_1273_), .B(_45_), .C(_47_), .Y(_48_) );
AND2X2 AND2X2_22 ( .A(_1221_), .B(_1409_), .Y(_49_) );
NAND3X1 NAND3X1_80 ( .A(_42_), .B(_48_), .C(_49_), .Y(_50_) );
NOR2X1 NOR2X1_118 ( .A(_50_), .B(_1429_), .Y(_51_) );
OAI21X1 OAI21X1_126 ( .A(_1425_), .B(_1426_), .C(_51_), .Y(_1438__3_) );
NAND3X1 NAND3X1_81 ( .A(_1117_), .B(_1152_), .C(_52_), .Y(_53_) );
AND2X2 AND2X2_23 ( .A(_1242_), .B(_1381_), .Y(_54_) );
NAND3X1 NAND3X1_82 ( .A(_1378_), .B(_54_), .C(_1434_), .Y(_55_) );
OR2X2 OR2X2_12 ( .A(_55_), .B(_53_), .Y(_56_) );
NOR2X1 NOR2X1_119 ( .A(_45_), .B(_56_), .Y(_57_) );
OAI21X1 OAI21X1_127 ( .A(new_wire_8), .B(_1320_), .C(_1322_), .Y(_58_) );
NOR2X1 NOR2X1_120 ( .A(_1414_), .B(_58_), .Y(_59_) );
NAND3X1 NAND3X1_83 ( .A(_1261_), .B(_1270_), .C(_1284_), .Y(_60_) );
NOR2X1 NOR2X1_121 ( .A(_1406_), .B(_60_), .Y(_61_) );
NAND3X1 NAND3X1_84 ( .A(_57_), .B(_59_), .C(_61_), .Y(_1438__4_) );
AND2X2 AND2X2_24 ( .A(_1239_), .B(_1238_), .Y(_62_) );
NOR2X1 NOR2X1_122 ( .A(_1314_), .B(_63_), .Y(_64_) );
NOR2X1 NOR2X1_123 ( .A(_1164_), .B(_65_), .Y(_66_) );
NOR2X1 NOR2X1_124 ( .A(_1121_), .B(_1113_), .Y(_67_) );
NOR2X1 NOR2X1_125 ( .A(_1204_), .B(_1157_), .Y(_68_) );
AND2X2 AND2X2_25 ( .A(_68_), .B(_67_), .Y(_69_) );
NAND3X1 NAND3X1_85 ( .A(_64_), .B(_66_), .C(_69_), .Y(_70_) );
AOI21X1 AOI21X1_49 ( .A(_1407_), .B(_1408_), .C(_71_), .Y(_72_) );
NAND3X1 NAND3X1_86 ( .A(_1142_), .B(_1383_), .C(_72_), .Y(_73_) );
NOR2X1 NOR2X1_126 ( .A(_73_), .B(_70_), .Y(_74_) );
NAND3X1 NAND3X1_87 ( .A(_62_), .B(_1411_), .C(_74_), .Y(_75_) );
NOR2X1 NOR2X1_127 ( .A(_1231_), .B(_1229_), .Y(_76_) );
NAND3X1 NAND3X1_88 ( .A(_1098_), .B(_1302_), .C(_76_), .Y(_77_) );
NOR2X1 NOR2X1_128 ( .A(_77_), .B(_75_), .Y(_78_) );
NAND3X1 NAND3X1_89 ( .A(_1391_), .B(_1393_), .C(_78_), .Y(_1438__5_) );
OAI21X1 OAI21X1_128 ( .A(_1196_), .B(_1210_), .C(new_wire_32), .Y(_80_) );
OAI21X1 OAI21X1_129 ( .A(_803_), .B(_809__bF_buf2), .C(_80_), .Y(_81_) );
OR2X2 OR2X2_13 ( .A(_1205_), .B(load_only), .Y(_82_) );
NOR2X1 NOR2X1_129 ( .A(shift), .B(_82_), .Y(_83_) );
AOI21X1 AOI21X1_50 ( .A(rotate), .B(_81_), .C(_83_), .Y(_84_) );
NAND3X1 NAND3X1_90 ( .A(inc), .B(_87_), .C(_88_), .Y(_89_) );
OAI21X1 OAI21X1_130 ( .A(_86_), .B(_1205_), .C(_89_), .Y(_90_) );
OAI21X1 OAI21X1_131 ( .A(_809__bF_buf3), .B(_1236_), .C(_815__bF_buf1), .Y(_92_) );
OAI21X1 OAI21X1_132 ( .A(_91_), .B(_92_), .C(CO), .Y(_93_) );
OAI21X1 OAI21X1_133 ( .A(_799__bF_buf4), .B(_1161_), .C(_1154_), .Y(_94_) );
OAI21X1 OAI21X1_134 ( .A(_799__bF_buf4), .B(_1171_), .C(_1230_), .Y(_95_) );
OR2X2 OR2X2_14 ( .A(_94_), .B(_95_), .Y(_96_) );
OAI21X1 OAI21X1_135 ( .A(_799__bF_buf3), .B(_792_), .C(_1143_), .Y(_98_) );
NAND3X1 NAND3X1_91 ( .A(_1320_), .B(_97_), .C(_99_), .Y(_100_) );
NOR2X1 NOR2X1_130 ( .A(_100_), .B(_96_), .Y(_101_) );
NAND2X1 NAND2X1_121 ( .A(_93_), .B(_101_), .Y(_102_) );
AOI21X1 AOI21X1_51 ( .A(_85_), .B(_90_), .C(_102_), .Y(_103_) );
OAI21X1 OAI21X1_136 ( .A(_79_), .B(_84_), .C(_103_), .Y(CI) );
NOR2X1 NOR2X1_131 ( .A(_1291_), .B(_88_), .Y(_105_) );
AOI21X1 AOI21X1_52 ( .A(_841_), .B(_812__bF_buf2), .C(_1170_), .Y(_106_) );
NOR2X1 NOR2X1_132 ( .A(_849__bF_buf4), .B(_1245_), .Y(_107_) );
NAND2X1 NAND2X1_122 ( .A(_107_), .B(_106_), .Y(_108_) );
NOR2X1 NOR2X1_133 ( .A(_840_), .B(_1195_), .Y(_109_) );
OAI21X1 OAI21X1_137 ( .A(_856_), .B(_109_), .C(_812__bF_buf1), .Y(_110_) );
NOR2X1 NOR2X1_134 ( .A(_1072_), .B(_1251_), .Y(_111_) );
NAND2X1 NAND2X1_123 ( .A(_110_), .B(_111_), .Y(_112_) );
NOR2X1 NOR2X1_135 ( .A(_108_), .B(_112_), .Y(_113_) );
NAND3X1 NAND3X1_92 ( .A(_114_), .B(_99_), .C(_1100_), .Y(_115_) );
NOR2X1 NOR2X1_136 ( .A(_96_), .B(_115_), .Y(_116_) );
NAND3X1 NAND3X1_93 ( .A(_105_), .B(_113_), .C(_116_), .Y(_117_) );
OAI22X1 OAI22X1_11 ( .A(_905_), .B(_1100_), .C(_104_), .D(_117_), .Y(BI_0_) );
OAI22X1 OAI22X1_12 ( .A(_933_), .B(_1100_), .C(_118_), .D(_117_), .Y(BI_1_) );
OAI22X1 OAI22X1_13 ( .A(_956_), .B(_1100_), .C(_978_), .D(_117_), .Y(BI_2_) );
OAI22X1 OAI22X1_14 ( .A(_944_), .B(_1100_), .C(_1179_), .D(_117_), .Y(BI_3_) );
OAI22X1 OAI22X1_15 ( .A(_872_), .B(_1100_), .C(_1019_), .D(_117_), .Y(BI_4_) );
OAI22X1 OAI22X1_16 ( .A(_860_), .B(new_wire_55), .C(_119_), .D(_117_), .Y(BI_5_) );
OAI22X1 OAI22X1_17 ( .A(_893_), .B(new_wire_55), .C(_1052_), .D(_117_), .Y(BI_6_) );
OAI22X1 OAI22X1_18 ( .A(_883_), .B(new_wire_55), .C(_1064_), .D(_117_), .Y(BI_7_) );
NOR2X1 NOR2X1_137 ( .A(_1006_), .B(_815__bF_buf3), .Y(_120_) );
OAI21X1 OAI21X1_138 ( .A(_809__bF_buf2), .B(_1171_), .C(_106_), .Y(_121_) );
OR2X2 OR2X2_15 ( .A(_121_), .B(_94_), .Y(_122_) );
OAI21X1 OAI21X1_139 ( .A(_98_), .B(_122_), .C(ADD_0_), .Y(_123_) );
OAI21X1 OAI21X1_140 ( .A(_799__bF_buf3), .B(_1236_), .C(new_wire_55), .Y(_124_) );
OAI21X1 OAI21X1_141 ( .A(_104_), .B(_125_), .C(_123_), .Y(_126_) );
NOR2X1 NOR2X1_138 ( .A(_120_), .B(_126_), .Y(_127_) );
OAI21X1 OAI21X1_142 ( .A(_809__bF_buf0), .B(_915_), .C(_1110_), .Y(_129_) );
OAI22X1 OAI22X1_19 ( .A(_795__bF_buf4), .B(_1236_), .C(_809__bF_buf3), .D(_1145_), .Y(_130_) );
NOR3X1 NOR3X1_12 ( .A(_859__bF_buf2), .B(_129_), .C(_130_), .Y(_131_) );
OAI22X1 OAI22X1_20 ( .A(_809__bF_buf2), .B(_1119_), .C(_795__bF_buf3), .D(_1171_), .Y(_132_) );
OAI21X1 OAI21X1_143 ( .A(_799__bF_buf3), .B(_1119_), .C(_1160_), .Y(_133_) );
NOR2X1 NOR2X1_139 ( .A(_132_), .B(_133_), .Y(_134_) );
OAI21X1 OAI21X1_144 ( .A(_795__bF_buf4), .B(_1145_), .C(_916_), .Y(_135_) );
NAND2X1 NAND2X1_124 ( .A(new_wire_31), .B(_1137_), .Y(_136_) );
OAI21X1 OAI21X1_145 ( .A(_799__bF_buf3), .B(_915_), .C(_136_), .Y(_137_) );
NAND3X1 NAND3X1_94 ( .A(_1201_), .B(_1244_), .C(_1230_), .Y(_138_) );
NOR3X1 NOR3X1_13 ( .A(_137_), .B(_135_), .C(_138_), .Y(_139_) );
NAND3X1 NAND3X1_95 ( .A(_131_), .B(_139_), .C(_134_), .Y(_140_) );
NOR2X1 NOR2X1_140 ( .A(_129_), .B(_130_), .Y(_142_) );
OAI21X1 OAI21X1_146 ( .A(_141_), .B(_822__bF_buf0), .C(_142_), .Y(_143_) );
OAI21X1 OAI21X1_147 ( .A(_128_), .B(_140_), .C(_144_), .Y(_145_) );
OR2X2 OR2X2_16 ( .A(_140_), .B(src_reg_0_), .Y(_148_) );
OAI21X1 OAI21X1_148 ( .A(_809__bF_buf3), .B(_811_), .C(_142_), .Y(_149_) );
OAI21X1 OAI21X1_149 ( .A(_129_), .B(_130_), .C(index_y), .Y(_150_) );
NAND2X1 NAND2X1_125 ( .A(dst_reg_0_), .B(_859__bF_buf2), .Y(_151_) );
NAND3X1 NAND3X1_96 ( .A(_150_), .B(_151_), .C(_149_), .Y(_152_) );
NAND3X1 NAND3X1_97 ( .A(_147_), .B(_152__bF_buf3), .C(_148__bF_buf2), .Y(_153_) );
OAI21X1 OAI21X1_150 ( .A(src_reg_0_), .B(_140_), .C(_152__bF_buf1), .Y(_155_) );
NAND2X1 NAND2X1_126 ( .A(_154_), .B(_155__bF_buf1), .Y(_156_) );
NAND3X1 NAND3X1_98 ( .A(_146_), .B(_156_), .C(_153_), .Y(_157_) );
NAND3X1 NAND3X1_99 ( .A(_158_), .B(_152__bF_buf3), .C(_148__bF_buf2), .Y(_159_) );
NAND2X1 NAND2X1_127 ( .A(_160_), .B(_155__bF_buf3), .Y(_161_) );
NAND3X1 NAND3X1_100 ( .A(_145_), .B(_161_), .C(_159_), .Y(_162_) );
AND2X2 AND2X2_26 ( .A(_157_), .B(_162_), .Y(_163_) );
NOR2X1 NOR2X1_141 ( .A(_1072_), .B(_1123_), .Y(_164_) );
OAI21X1 OAI21X1_151 ( .A(_920_), .B(_1319_), .C(new_wire_32), .Y(_165_) );
OAI21X1 OAI21X1_152 ( .A(new_wire_31), .B(new_wire_32), .C(_856_), .Y(_166_) );
AND2X2 AND2X2_27 ( .A(_165_), .B(_166_), .Y(_167_) );
NAND3X1 NAND3X1_101 ( .A(_82_), .B(_164_), .C(_167_), .Y(_168_) );
NOR2X1 NOR2X1_142 ( .A(_1245_), .B(_1251_), .Y(_170_) );
NAND3X1 NAND3X1_102 ( .A(_169_), .B(_170_), .C(_142_), .Y(_171_) );
NOR2X1 NOR2X1_143 ( .A(_171_), .B(_168_), .Y(_172_) );
OAI21X1 OAI21X1_153 ( .A(_172_), .B(_163_), .C(_127_), .Y(AI_0_) );
OR2X2 OR2X2_17 ( .A(_122_), .B(_98_), .Y(_173_) );
OAI22X1 OAI22X1_21 ( .A(_994_), .B(_815__bF_buf3), .C(_118_), .D(_125_), .Y(_174_) );
AOI21X1 AOI21X1_53 ( .A(_173_), .B(ADD_1_), .C(_174_), .Y(_175_) );
NAND3X1 NAND3X1_103 ( .A(_176_), .B(_152__bF_buf1), .C(_148__bF_buf0), .Y(_177_) );
NAND2X1 NAND2X1_128 ( .A(_178_), .B(_155__bF_buf0), .Y(_179_) );
NAND3X1 NAND3X1_104 ( .A(_146_), .B(_179_), .C(_177_), .Y(_180_) );
NAND3X1 NAND3X1_105 ( .A(_181_), .B(_152__bF_buf3), .C(_148__bF_buf0), .Y(_182_) );
NAND2X1 NAND2X1_129 ( .A(_183_), .B(_155__bF_buf3), .Y(_184_) );
NAND3X1 NAND3X1_106 ( .A(_145_), .B(_184_), .C(_182_), .Y(_185_) );
AND2X2 AND2X2_28 ( .A(_180_), .B(_185_), .Y(_186_) );
OAI21X1 OAI21X1_154 ( .A(_172_), .B(_186_), .C(_175_), .Y(AI_1_) );
OAI22X1 OAI22X1_22 ( .A(_981_), .B(_815__bF_buf3), .C(_978_), .D(_125_), .Y(_187_) );
AOI21X1 AOI21X1_54 ( .A(_173_), .B(ADD_2_), .C(_187_), .Y(_188_) );
NAND3X1 NAND3X1_107 ( .A(_189_), .B(_152__bF_buf2), .C(_148__bF_buf3), .Y(_190_) );
NAND2X1 NAND2X1_130 ( .A(_191_), .B(_155__bF_buf2), .Y(_192_) );
NAND3X1 NAND3X1_108 ( .A(_146_), .B(_192_), .C(_190_), .Y(_193_) );
NAND3X1 NAND3X1_109 ( .A(_194_), .B(_152__bF_buf2), .C(_148__bF_buf3), .Y(_195_) );
NAND2X1 NAND2X1_131 ( .A(_196_), .B(_155__bF_buf2), .Y(_197_) );
NAND3X1 NAND3X1_110 ( .A(_145_), .B(_197_), .C(_195_), .Y(_198_) );
AND2X2 AND2X2_29 ( .A(_193_), .B(_198_), .Y(_199_) );
OAI21X1 OAI21X1_155 ( .A(_172_), .B(_199_), .C(_188_), .Y(AI_2_) );
OAI22X1 OAI22X1_23 ( .A(_970_), .B(_815__bF_buf3), .C(_1179_), .D(_125_), .Y(_200_) );
AOI21X1 AOI21X1_55 ( .A(_173_), .B(ADD_3_), .C(_200_), .Y(_201_) );
NAND3X1 NAND3X1_111 ( .A(_202_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_203_) );
NAND2X1 NAND2X1_132 ( .A(_204_), .B(_155__bF_buf3), .Y(_205_) );
NAND3X1 NAND3X1_112 ( .A(_146_), .B(_205_), .C(_203_), .Y(_206_) );
NAND3X1 NAND3X1_113 ( .A(_207_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_208_) );
NAND2X1 NAND2X1_133 ( .A(_209_), .B(_155__bF_buf0), .Y(_210_) );
NAND3X1 NAND3X1_114 ( .A(_145_), .B(_210_), .C(_208_), .Y(_211_) );
AND2X2 AND2X2_30 ( .A(_206_), .B(_211_), .Y(_212_) );
OAI21X1 OAI21X1_156 ( .A(_172_), .B(_212_), .C(_201_), .Y(AI_3_) );
OAI22X1 OAI22X1_24 ( .A(_1020_), .B(_815__bF_buf3), .C(_1019_), .D(_125_), .Y(_213_) );
AOI21X1 AOI21X1_56 ( .A(_173_), .B(ADD_4_), .C(_213_), .Y(_214_) );
NAND3X1 NAND3X1_115 ( .A(_215_), .B(_152__bF_buf1), .C(_148__bF_buf0), .Y(_216_) );
NAND2X1 NAND2X1_134 ( .A(_217_), .B(_155__bF_buf0), .Y(_218_) );
NAND3X1 NAND3X1_116 ( .A(_146_), .B(_218_), .C(_216_), .Y(_219_) );
NAND3X1 NAND3X1_117 ( .A(_220_), .B(_152__bF_buf1), .C(_148__bF_buf0), .Y(_221_) );
NAND2X1 NAND2X1_135 ( .A(_222_), .B(_155__bF_buf3), .Y(_223_) );
NAND3X1 NAND3X1_118 ( .A(_145_), .B(_223_), .C(_221_), .Y(_224_) );
AND2X2 AND2X2_31 ( .A(_219_), .B(_224_), .Y(_225_) );
OAI21X1 OAI21X1_157 ( .A(_172_), .B(_225_), .C(_214_), .Y(AI_4_) );
OAI22X1 OAI22X1_25 ( .A(_226_), .B(_815__bF_buf2), .C(_119_), .D(_125_), .Y(_227_) );
AOI21X1 AOI21X1_57 ( .A(_173_), .B(ADD_5_), .C(_227_), .Y(_228_) );
NAND3X1 NAND3X1_119 ( .A(_229_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_230_) );
NAND2X1 NAND2X1_136 ( .A(_231_), .B(_155__bF_buf1), .Y(_232_) );
NAND3X1 NAND3X1_120 ( .A(_146_), .B(_232_), .C(_230_), .Y(_233_) );
NAND3X1 NAND3X1_121 ( .A(_234_), .B(_152__bF_buf0), .C(_148__bF_buf1), .Y(_235_) );
NAND2X1 NAND2X1_137 ( .A(_236_), .B(_155__bF_buf3), .Y(_237_) );
NAND3X1 NAND3X1_122 ( .A(_145_), .B(_237_), .C(_235_), .Y(_238_) );
AND2X2 AND2X2_32 ( .A(_233_), .B(_238_), .Y(_239_) );
OAI21X1 OAI21X1_158 ( .A(_172_), .B(_239_), .C(_228_), .Y(AI_5_) );
OAI22X1 OAI22X1_26 ( .A(_1049_), .B(_815__bF_buf2), .C(_1052_), .D(_125_), .Y(_240_) );
AOI21X1 AOI21X1_58 ( .A(_173_), .B(ADD_6_), .C(_240_), .Y(_241_) );
NAND3X1 NAND3X1_123 ( .A(_242_), .B(_152__bF_buf3), .C(_148__bF_buf2), .Y(_243_) );
NAND2X1 NAND2X1_138 ( .A(_244_), .B(_155__bF_buf1), .Y(_245_) );
NAND3X1 NAND3X1_124 ( .A(_146_), .B(_245_), .C(_243_), .Y(_246_) );
NAND3X1 NAND3X1_125 ( .A(_247_), .B(_152__bF_buf3), .C(_148__bF_buf2), .Y(_248_) );
NAND2X1 NAND2X1_139 ( .A(_249_), .B(_155__bF_buf1), .Y(_250_) );
NAND3X1 NAND3X1_126 ( .A(_145_), .B(_250_), .C(_248_), .Y(_251_) );
AND2X2 AND2X2_33 ( .A(_246_), .B(_251_), .Y(_252_) );
OAI21X1 OAI21X1_159 ( .A(_172_), .B(_252_), .C(_241_), .Y(AI_6_) );
OAI22X1 OAI22X1_27 ( .A(_1061_), .B(_815__bF_buf2), .C(_1064_), .D(_125_), .Y(_253_) );
AOI21X1 AOI21X1_59 ( .A(_173_), .B(ADD_7_), .C(_253_), .Y(_254_) );
NAND3X1 NAND3X1_127 ( .A(_255_), .B(_152__bF_buf2), .C(_148__bF_buf3), .Y(_256_) );
NAND2X1 NAND2X1_140 ( .A(_257_), .B(_155__bF_buf2), .Y(_258_) );
NAND3X1 NAND3X1_128 ( .A(_146_), .B(_258_), .C(_256_), .Y(_259_) );
NAND3X1 NAND3X1_129 ( .A(_260_), .B(_152__bF_buf2), .C(_148__bF_buf3), .Y(_261_) );
NAND2X1 NAND2X1_141 ( .A(_262_), .B(_155__bF_buf2), .Y(_263_) );
NAND3X1 NAND3X1_130 ( .A(new_wire_61), .B(_263_), .C(_261_), .Y(_264_) );
AND2X2 AND2X2_34 ( .A(_259_), .B(_264_), .Y(_265_) );
OAI21X1 OAI21X1_160 ( .A(_172_), .B(_265_), .C(_254_), .Y(AI_7_) );
NOR3X1 NOR3X1_14 ( .A(_816_), .B(_1130_), .C(_81_), .Y(_268_) );
OAI21X1 OAI21X1_161 ( .A(_799__bF_buf4), .B(_915_), .C(_269_), .Y(_270_) );
NOR2X1 NOR2X1_144 ( .A(_270_), .B(_121_), .Y(_271_) );
NAND2X1 NAND2X1_142 ( .A(_815__bF_buf2), .B(_271_), .Y(_272_) );
NOR2X1 NOR2X1_145 ( .A(_268_), .B(_272_), .Y(_273_) );
OAI21X1 OAI21X1_162 ( .A(_266_), .B(_267_), .C(_273_), .Y(alu_op_0_) );
OAI21X1 OAI21X1_163 ( .A(_274_), .B(_267_), .C(_273_), .Y(alu_op_1_) );
AOI21X1 AOI21X1_60 ( .A(op_2_), .B(_81_), .C(_276_), .Y(_277_) );
OAI21X1 OAI21X1_164 ( .A(_275_), .B(_815__bF_buf1), .C(_277_), .Y(alu_op_2_) );
NOR2X1 NOR2X1_146 ( .A(_278_), .B(_267_), .Y(alu_op_3_) );
OAI21X1 OAI21X1_165 ( .A(_799__bF_buf3), .B(_1145_), .C(_271_), .Y(_280_) );
AND2X2 AND2X2_35 ( .A(_1199_), .B(_1190_), .Y(_282_) );
OAI21X1 OAI21X1_166 ( .A(_279_), .B(_282_), .C(_281_), .Y(_1441_) );
MUX2X1 MUX2X1_10 ( .A(C), .B(ADD_0_), .S(php), .Y(_284_) );
OAI22X1 OAI22X1_28 ( .A(_79_), .B(_817_), .C(_284_), .D(_114_), .Y(_285_) );
AOI21X1 AOI21X1_61 ( .A(ADD_0_), .B(_283_), .C(_285_), .Y(_286_) );
AOI22X1 AOI22X1_26 ( .A(PC_8_), .B(_132_), .C(PC_0_), .D(_287_), .Y(_288_) );
AND2X2 AND2X2_36 ( .A(_286_), .B(_288_), .Y(_289_) );
OAI21X1 OAI21X1_167 ( .A(_280_), .B(_163_), .C(_289_), .Y(_1440__0_) );
OAI21X1 OAI21X1_168 ( .A(_290_), .B(_114_), .C(_817_), .Y(_291_) );
AOI22X1 AOI22X1_27 ( .A(PC_9_), .B(_132_), .C(PC_1_), .D(_287_), .Y(_292_) );
OAI21X1 OAI21X1_169 ( .A(php), .B(_114_), .C(_1192_), .Y(_293_) );
OAI21X1 OAI21X1_170 ( .A(_931_), .B(_294_), .C(_292_), .Y(_295_) );
AOI21X1 AOI21X1_62 ( .A(Z), .B(_291_), .C(_295_), .Y(_296_) );
OAI21X1 OAI21X1_171 ( .A(_280_), .B(_186_), .C(_296_), .Y(_1440__1_) );
NAND2X1 NAND2X1_143 ( .A(ADD_2_), .B(_293_), .Y(_297_) );
OAI22X1 OAI22X1_29 ( .A(_983_), .B(_269_), .C(_956_), .D(_106_), .Y(_298_) );
AOI21X1 AOI21X1_63 ( .A(I), .B(_291_), .C(_298_), .Y(_299_) );
AND2X2 AND2X2_37 ( .A(_299_), .B(_297_), .Y(_300_) );
OAI21X1 OAI21X1_172 ( .A(_280_), .B(_199_), .C(_300_), .Y(_1440__2_) );
NOR2X1 NOR2X1_147 ( .A(_290_), .B(_114_), .Y(_301_) );
OAI21X1 OAI21X1_173 ( .A(new_wire_43), .B(_301_), .C(D), .Y(_302_) );
OAI22X1 OAI22X1_30 ( .A(_972_), .B(_269_), .C(_944_), .D(_106_), .Y(_303_) );
AOI21X1 AOI21X1_64 ( .A(ADD_3_), .B(_293_), .C(_303_), .Y(_304_) );
AND2X2 AND2X2_38 ( .A(_304_), .B(_302_), .Y(_305_) );
OAI21X1 OAI21X1_174 ( .A(_280_), .B(_212_), .C(_305_), .Y(_1440__3_) );
OAI22X1 OAI22X1_31 ( .A(_283_), .B(_1323_), .C(ADD_4_), .D(_301_), .Y(_306_) );
OAI21X1 OAI21X1_175 ( .A(new_wire_34), .B(_829_), .C(_306_), .Y(_307_) );
OAI22X1 OAI22X1_32 ( .A(_1016_), .B(_269_), .C(_872_), .D(_106_), .Y(_308_) );
NOR2X1 NOR2X1_148 ( .A(_308_), .B(_307_), .Y(_309_) );
OAI21X1 OAI21X1_176 ( .A(_280_), .B(_225_), .C(_309_), .Y(_1440__4_) );
OAI22X1 OAI22X1_33 ( .A(_283_), .B(_1323_), .C(ADD_5_), .D(_301_), .Y(_310_) );
OAI21X1 OAI21X1_177 ( .A(_787_), .B(_269_), .C(new_wire_34), .Y(_311_) );
AOI21X1 AOI21X1_65 ( .A(PC_5_), .B(_287_), .C(_311_), .Y(_312_) );
AND2X2 AND2X2_39 ( .A(_312_), .B(_310_), .Y(_313_) );
OAI21X1 OAI21X1_178 ( .A(_280_), .B(_239_), .C(_313_), .Y(_1440__5_) );
AOI22X1 AOI22X1_28 ( .A(PC_14_), .B(_132_), .C(PC_6_), .D(_287_), .Y(_315_) );
OAI21X1 OAI21X1_179 ( .A(_1306_), .B(_314_), .C(_315_), .Y(_316_) );
AOI21X1 AOI21X1_66 ( .A(ADD_6_), .B(_293_), .C(_316_), .Y(_317_) );
OAI21X1 OAI21X1_180 ( .A(_280_), .B(_252_), .C(_317_), .Y(_1440__6_) );
AOI22X1 AOI22X1_29 ( .A(PC_15_), .B(_132_), .C(PC_7_), .D(_287_), .Y(_319_) );
OAI21X1 OAI21X1_181 ( .A(_318_), .B(_314_), .C(_319_), .Y(_320_) );
AOI21X1 AOI21X1_67 ( .A(ADD_7_), .B(_293_), .C(_320_), .Y(_321_) );
OAI21X1 OAI21X1_182 ( .A(new_wire_67), .B(_265_), .C(_321_), .Y(_1440__7_) );
AND2X2 AND2X2_40 ( .A(D), .B(adc_sbc), .Y(_14_) );
NOR2X1 NOR2X1_149 ( .A(_322_), .B(_1205_), .Y(ALU_BCD) );
OAI21X1 OAI21X1_183 ( .A(_323_), .B(_859__bF_buf0), .C(_1175_), .Y(_31_) );
NOR2X1 NOR2X1_150 ( .A(_324_), .B(_822__bF_buf2), .Y(_325_) );
OAI21X1 OAI21X1_184 ( .A(_828_), .B(_325_), .C(_169_), .Y(_326_) );
AOI21X1 AOI21X1_68 ( .A(ADD_2_), .B(_325_), .C(_326_), .Y(_327_) );
AOI21X1 AOI21X1_69 ( .A(_1155_), .B(DIMUX_2_), .C(_328_), .Y(_329_) );
AOI21X1 AOI21X1_70 ( .A(_828_), .B(_331_), .C(cli), .Y(_332_) );
OAI21X1 OAI21X1_185 ( .A(_332_), .B(_169_), .C(_330_), .Y(_333_) );
OAI21X1 OAI21X1_186 ( .A(_333_), .B(_327_), .C(_329_), .Y(_6_) );
AND2X2 AND2X2_41 ( .A(_81_), .B(shift_right), .Y(alu_shift_right) );
OAI21X1 OAI21X1_187 ( .A(_811_), .B(_795__bF_buf3), .C(_916_), .Y(_334_) );
OAI21X1 OAI21X1_188 ( .A(_795__bF_buf3), .B(_1171_), .C(_136_), .Y(_335_) );
NOR2X1 NOR2X1_151 ( .A(_334_), .B(_335_), .Y(_336_) );
OAI21X1 OAI21X1_189 ( .A(_799__bF_buf4), .B(_1119_), .C(_1201_), .Y(_337_) );
NOR2X1 NOR2X1_152 ( .A(plp), .B(_338_), .Y(_339_) );
AOI21X1 AOI21X1_71 ( .A(_859__bF_buf2), .B(_339_), .C(_337_), .Y(_340_) );
AOI21X1 AOI21X1_72 ( .A(_336_), .B(_340_), .C(_1017__bF_buf2), .Y(_341_) );
NAND3X1 NAND3X1_131 ( .A(_152__bF_buf2), .B(_341_), .C(_148__bF_buf3), .Y(_342_) );
NOR2X1 NOR2X1_153 ( .A(new_wire_61), .B(_342_), .Y(_343_) );
OAI21X1 OAI21X1_190 ( .A(_795__bF_buf3), .B(_1171_), .C(_904_), .Y(_344_) );
OAI21X1 OAI21X1_191 ( .A(DIMUX_0_), .B(_43_), .C(_344_), .Y(_345_) );
MUX2X1 MUX2X1_11 ( .A(_345_), .B(_147_), .S(_343_), .Y(_1442__0_) );
NOR2X1 NOR2X1_154 ( .A(adc_bcd), .B(HC), .Y(_346_) );
NAND2X1 NAND2X1_144 ( .A(adj_bcd), .B(_346_), .Y(_347_) );
NAND3X1 NAND3X1_132 ( .A(adc_bcd), .B(adj_bcd), .C(HC), .Y(_348_) );
NAND2X1 NAND2X1_145 ( .A(_348_), .B(_347_), .Y(_349_) );
NAND2X1 NAND2X1_146 ( .A(_931_), .B(_350_), .Y(_351_) );
NOR2X1 NOR2X1_155 ( .A(_931_), .B(_350_), .Y(_352_) );
NOR2X1 NOR2X1_156 ( .A(_1291_), .B(_352_), .Y(_353_) );
AOI22X1 AOI22X1_30 ( .A(DIMUX_1_), .B(_1291_), .C(_351_), .D(_353_), .Y(_354_) );
MUX2X1 MUX2X1_12 ( .A(_354_), .B(_176_), .S(_343_), .Y(_1442__1_) );
XNOR2X1 XNOR2X1_2 ( .A(_348_), .B(ADD_2_), .Y(_355_) );
OAI21X1 OAI21X1_192 ( .A(_931_), .B(_350_), .C(_356_), .Y(_357_) );
AOI21X1 AOI21X1_73 ( .A(_352_), .B(_355_), .C(_1291_), .Y(_358_) );
AOI22X1 AOI22X1_31 ( .A(DIMUX_2_), .B(_1291_), .C(_357_), .D(_358_), .Y(_359_) );
MUX2X1 MUX2X1_13 ( .A(_359_), .B(_189_), .S(_343_), .Y(_1442__2_) );
NAND2X1 NAND2X1_147 ( .A(_355_), .B(_352_), .Y(_361_) );
OAI21X1 OAI21X1_193 ( .A(_360_), .B(_348_), .C(_361_), .Y(_362_) );
XNOR2X1 XNOR2X1_3 ( .A(_347_), .B(_363_), .Y(_364_) );
XNOR2X1 XNOR2X1_4 ( .A(_362_), .B(_364_), .Y(_365_) );
MUX2X1 MUX2X1_14 ( .A(_365_), .B(DIMUX_3_), .S(_43_), .Y(_366_) );
MUX2X1 MUX2X1_15 ( .A(_366_), .B(_202_), .S(_343_), .Y(_1442__3_) );
OAI21X1 OAI21X1_194 ( .A(_795__bF_buf3), .B(_1171_), .C(_367_), .Y(_368_) );
OAI21X1 OAI21X1_195 ( .A(DIMUX_4_), .B(_43_), .C(_368_), .Y(_369_) );
MUX2X1 MUX2X1_16 ( .A(_369_), .B(_215_), .S(_343_), .Y(_1442__4_) );
NAND3X1 NAND3X1_133 ( .A(adj_bcd), .B(_370_), .C(_322_), .Y(_371_) );
NAND3X1 NAND3X1_134 ( .A(CO), .B(adc_bcd), .C(adj_bcd), .Y(_372_) );
NAND2X1 NAND2X1_148 ( .A(_372_), .B(_371_), .Y(_373_) );
NAND2X1 NAND2X1_149 ( .A(_846_), .B(_374_), .Y(_375_) );
NOR2X1 NOR2X1_157 ( .A(_846_), .B(_374_), .Y(_376_) );
NOR2X1 NOR2X1_158 ( .A(_1291_), .B(_376_), .Y(_377_) );
AOI22X1 AOI22X1_32 ( .A(DIMUX_5_), .B(new_wire_59), .C(_375_), .D(_377_), .Y(_378_) );
MUX2X1 MUX2X1_17 ( .A(_378_), .B(_229_), .S(_343_), .Y(_1442__5_) );
XNOR2X1 XNOR2X1_5 ( .A(_372_), .B(ADD_6_), .Y(_379_) );
OAI21X1 OAI21X1_196 ( .A(_846_), .B(_374_), .C(_380_), .Y(_381_) );
AOI21X1 AOI21X1_74 ( .A(_376_), .B(_379_), .C(new_wire_59), .Y(_382_) );
AOI22X1 AOI22X1_33 ( .A(DIMUX_6_), .B(new_wire_59), .C(_381_), .D(_382_), .Y(_383_) );
MUX2X1 MUX2X1_18 ( .A(_383_), .B(_242_), .S(_343_), .Y(_1442__6_) );
NAND2X1 NAND2X1_150 ( .A(_379_), .B(_376_), .Y(_385_) );
OAI21X1 OAI21X1_197 ( .A(_384_), .B(_372_), .C(_385_), .Y(_386_) );
XNOR2X1 XNOR2X1_6 ( .A(_371_), .B(_387_), .Y(_388_) );
XNOR2X1 XNOR2X1_7 ( .A(_386_), .B(_388_), .Y(_389_) );
MUX2X1 MUX2X1_19 ( .A(_389_), .B(DIMUX_7_), .S(_43_), .Y(_390_) );
MUX2X1 MUX2X1_20 ( .A(_390_), .B(_255_), .S(_343_), .Y(_1442__7_) );
NAND3X1 NAND3X1_135 ( .A(NMI), .B(new_wire_40), .C(_391_), .Y(_392_) );
OAI21X1 OAI21X1_198 ( .A(new_wire_40), .B(_328_), .C(_392_), .Y(_7_) );
NAND2X1 NAND2X1_151 ( .A(cond_code_0_), .B(_1017__bF_buf3), .Y(_393_) );
OAI21X1 OAI21X1_199 ( .A(_1017__bF_buf3), .B(_1361_), .C(_393_), .Y(_22__0_) );
NAND2X1 NAND2X1_152 ( .A(cond_code_1_), .B(_1017__bF_buf7), .Y(_394_) );
OAI21X1 OAI21X1_200 ( .A(_1017__bF_buf7), .B(_1226_), .C(_394_), .Y(_22__1_) );
NAND2X1 NAND2X1_153 ( .A(cond_code_2_), .B(_1017__bF_buf7), .Y(_395_) );
OAI21X1 OAI21X1_201 ( .A(new_wire_22), .B(_1090_), .C(_395_), .Y(_22__2_) );
NAND2X1 NAND2X1_154 ( .A(_1070__bF_buf0), .B(_1266_), .Y(_396_) );
OAI22X1 OAI22X1_34 ( .A(_324_), .B(_1070__bF_buf2), .C(_1294_), .D(_396_), .Y(_30_) );
NOR2X1 NOR2X1_159 ( .A(_1101__bF_buf1), .B(_1275_), .Y(_398_) );
OAI22X1 OAI22X1_35 ( .A(_290_), .B(_1070__bF_buf2), .C(_399_), .D(_397_), .Y(_29_) );
OAI21X1 OAI21X1_202 ( .A(_1017__bF_buf3), .B(_822__bF_buf1), .C(clc), .Y(_400_) );
OAI21X1 OAI21X1_203 ( .A(_825__bF_buf0), .B(_1093_), .C(new_wire_56), .Y(_401_) );
NAND3X1 NAND3X1_136 ( .A(_1090_), .B(_398_), .C(_1266_), .Y(_402_) );
OAI21X1 OAI21X1_204 ( .A(_401_), .B(_402_), .C(_400_), .Y(_17_) );
OAI21X1 OAI21X1_205 ( .A(_1017__bF_buf1), .B(_822__bF_buf4), .C(sec), .Y(_403_) );
NOR2X1 NOR2X1_160 ( .A(new_wire_58), .B(_1361_), .Y(_404_) );
OAI21X1 OAI21X1_206 ( .A(_405_), .B(_402_), .C(_403_), .Y(_33_) );
OAI21X1 OAI21X1_207 ( .A(_1017__bF_buf3), .B(_822__bF_buf1), .C(cld), .Y(_406_) );
OR2X2 OR2X2_18 ( .A(_401_), .B(_1101__bF_buf0), .Y(_407_) );
NOR2X1 NOR2X1_161 ( .A(_1090_), .B(_1226_), .Y(_408_) );
NAND2X1 NAND2X1_155 ( .A(_408_), .B(_1266_), .Y(_409_) );
OAI21X1 OAI21X1_208 ( .A(_407_), .B(_409_), .C(_406_), .Y(_18_) );
OAI21X1 OAI21X1_209 ( .A(_1017__bF_buf3), .B(_822__bF_buf1), .C(sed), .Y(_410_) );
NAND2X1 NAND2X1_156 ( .A(_1070__bF_buf0), .B(_404_), .Y(_411_) );
OAI21X1 OAI21X1_210 ( .A(_411_), .B(_409_), .C(_410_), .Y(_34_) );
OAI21X1 OAI21X1_211 ( .A(_1017__bF_buf1), .B(_822__bF_buf1), .C(cli), .Y(_412_) );
NOR2X1 NOR2X1_162 ( .A(_1226_), .B(_1267_), .Y(_413_) );
NAND2X1 NAND2X1_157 ( .A(_413_), .B(_1266_), .Y(_414_) );
OAI21X1 OAI21X1_212 ( .A(_407_), .B(_414_), .C(_412_), .Y(_19_) );
OAI22X1 OAI22X1_36 ( .A(_331_), .B(_1070__bF_buf0), .C(_411_), .D(_414_), .Y(_35_) );
NOR2X1 NOR2X1_163 ( .A(_1090_), .B(_1275_), .Y(_415_) );
NAND2X1 NAND2X1_158 ( .A(_415_), .B(_404_), .Y(_416_) );
OAI21X1 OAI21X1_213 ( .A(_1017__bF_buf3), .B(_822__bF_buf0), .C(clv), .Y(_417_) );
OAI21X1 OAI21X1_214 ( .A(_416_), .B(_396_), .C(_417_), .Y(_20_) );
OAI21X1 OAI21X1_215 ( .A(_825__bF_buf3), .B(_1084_), .C(_1080_), .Y(_418_) );
OAI21X1 OAI21X1_216 ( .A(_825__bF_buf0), .B(_1082_), .C(_419_), .Y(_420_) );
OR2X2 OR2X2_19 ( .A(_420_), .B(_1294_), .Y(_421_) );
OAI21X1 OAI21X1_217 ( .A(_1017__bF_buf1), .B(_822__bF_buf4), .C(bit_ins), .Y(_422_) );
OAI21X1 OAI21X1_218 ( .A(_1101__bF_buf2), .B(_421_), .C(_422_), .Y(_16_) );
NAND2X1 NAND2X1_159 ( .A(new_wire_53), .B(_1388_), .Y(_423_) );
NOR2X1 NOR2X1_164 ( .A(_1140_), .B(_1094_), .Y(_426_) );
AOI21X1 AOI21X1_75 ( .A(_1388_), .B(_426_), .C(_425_), .Y(_427_) );
NAND3X1 NAND3X1_137 ( .A(_1267_), .B(_1095_), .C(_1266_), .Y(_428_) );
OAI22X1 OAI22X1_37 ( .A(_424_), .B(_427_), .C(_1275_), .D(_428_), .Y(_429_) );
NOR2X1 NOR2X1_165 ( .A(_1265_), .B(_424_), .Y(_430_) );
NOR2X1 NOR2X1_166 ( .A(new_wire_56), .B(_424_), .Y(_431_) );
AOI22X1 AOI22X1_34 ( .A(_430_), .B(_1136_), .C(_1279_), .D(_431_), .Y(_432_) );
NAND3X1 NAND3X1_138 ( .A(_1187_), .B(_1227_), .C(_1359_), .Y(_433_) );
NAND2X1 NAND2X1_160 ( .A(_433_), .B(_432_), .Y(_434_) );
NOR2X1 NOR2X1_167 ( .A(_429_), .B(_434_), .Y(_435_) );
NAND3X1 NAND3X1_139 ( .A(new_wire_53), .B(_1299_), .C(_425_), .Y(_436_) );
NAND2X1 NAND2X1_161 ( .A(_413_), .B(_1388_), .Y(_438_) );
OAI21X1 OAI21X1_219 ( .A(_1294_), .B(_420_), .C(_438_), .Y(_439_) );
NOR2X1 NOR2X1_168 ( .A(_437_), .B(_439_), .Y(_440_) );
NAND2X1 NAND2X1_162 ( .A(_440_), .B(_435_), .Y(_441_) );
OAI21X1 OAI21X1_220 ( .A(_1275_), .B(_423_), .C(_442_), .Y(_443_) );
NOR2X1 NOR2X1_169 ( .A(_1294_), .B(_420_), .Y(_445_) );
OAI21X1 OAI21X1_221 ( .A(_1267_), .B(_1358_), .C(_1070__bF_buf1), .Y(_446_) );
NOR2X1 NOR2X1_170 ( .A(_446_), .B(_445_), .Y(_447_) );
OAI21X1 OAI21X1_222 ( .A(_1361_), .B(_436_), .C(_447_), .Y(_448_) );
NOR2X1 NOR2X1_171 ( .A(_448_), .B(_444_), .Y(_449_) );
AOI22X1 AOI22X1_35 ( .A(_266_), .B(_1101__bF_buf2), .C(_449_), .D(_443_), .Y(_28__0_) );
NOR2X1 NOR2X1_172 ( .A(_1276_), .B(_1183_), .Y(_450_) );
AOI21X1 AOI21X1_76 ( .A(_450_), .B(new_wire_53), .C(_446_), .Y(_451_) );
AND2X2 AND2X2_42 ( .A(_435_), .B(_451_), .Y(_452_) );
AOI22X1 AOI22X1_36 ( .A(_274_), .B(_1101__bF_buf2), .C(_441_), .D(_452_), .Y(_28__1_) );
OAI21X1 OAI21X1_223 ( .A(_1017__bF_buf1), .B(_822__bF_buf4), .C(op_2_), .Y(_453_) );
OAI21X1 OAI21X1_224 ( .A(_1101__bF_buf2), .B(_442_), .C(_453_), .Y(_28__2_) );
AOI22X1 AOI22X1_37 ( .A(_278_), .B(_1101__bF_buf2), .C(_436_), .D(_447_), .Y(_28__3_) );
NAND3X1 NAND3X1_140 ( .A(_1083_), .B(_1094_), .C(_419_), .Y(_454_) );
NOR2X1 NOR2X1_173 ( .A(_1267_), .B(_454_), .Y(_455_) );
AOI21X1 AOI21X1_77 ( .A(_1362_), .B(_1359_), .C(_455_), .Y(_456_) );
OAI21X1 OAI21X1_225 ( .A(_1017__bF_buf1), .B(_822__bF_buf0), .C(rotate), .Y(_457_) );
OAI21X1 OAI21X1_226 ( .A(_1101__bF_buf0), .B(_456_), .C(_457_), .Y(_32_) );
OAI21X1 OAI21X1_227 ( .A(_1017__bF_buf1), .B(_822__bF_buf4), .C(shift_right), .Y(_458_) );
OAI21X1 OAI21X1_228 ( .A(_1101__bF_buf2), .B(_438_), .C(_458_), .Y(_37_) );
AOI21X1 AOI21X1_78 ( .A(_450_), .B(_1267_), .C(_1101__bF_buf0), .Y(_459_) );
AOI22X1 AOI22X1_38 ( .A(_86_), .B(_1101__bF_buf0), .C(_459_), .D(_432_), .Y(_21_) );
OAI21X1 OAI21X1_229 ( .A(_1080_), .B(_1181_), .C(_1070__bF_buf1), .Y(_460_) );
OAI22X1 OAI22X1_38 ( .A(_87_), .B(_1070__bF_buf0), .C(_460_), .D(_423_), .Y(_36_) );
OAI21X1 OAI21X1_230 ( .A(_859__bF_buf2), .B(_1123_), .C(RDY_bF_buf0), .Y(_461_) );
NAND2X1 NAND2X1_163 ( .A(D), .B(new_wire_53), .Y(_463_) );
NOR2X1 NOR2X1_174 ( .A(_1299_), .B(_1183_), .Y(_464_) );
NAND2X1 NAND2X1_164 ( .A(_462_), .B(_464_), .Y(_465_) );
OAI22X1 OAI22X1_39 ( .A(_322_), .B(_462_), .C(_463_), .D(_465_), .Y(_12_) );
OAI21X1 OAI21X1_231 ( .A(_466_), .B(_462_), .C(_465_), .Y(_13_) );
OAI21X1 OAI21X1_232 ( .A(new_wire_56), .B(_1087_), .C(_454_), .Y(_467_) );
NAND2X1 NAND2X1_165 ( .A(_408_), .B(_467_), .Y(_468_) );
OAI21X1 OAI21X1_233 ( .A(_1017__bF_buf1), .B(_822__bF_buf0), .C(inc), .Y(_469_) );
OAI21X1 OAI21X1_234 ( .A(_1101__bF_buf0), .B(_468_), .C(_469_), .Y(_24_) );
AND2X2 AND2X2_43 ( .A(_155__bF_buf2), .B(_341_), .Y(_470_) );
NAND2X1 NAND2X1_166 ( .A(new_wire_62), .B(_470_), .Y(_471_) );
NAND2X1 NAND2X1_167 ( .A(AXYS_0__0_), .B(_471_), .Y(_472_) );
OAI21X1 OAI21X1_235 ( .A(_345_), .B(_471_), .C(_472_), .Y(_1443__0_) );
NAND2X1 NAND2X1_168 ( .A(AXYS_0__1_), .B(_471_), .Y(_473_) );
OAI21X1 OAI21X1_236 ( .A(_354_), .B(_471_), .C(_473_), .Y(_1443__1_) );
NAND2X1 NAND2X1_169 ( .A(AXYS_0__2_), .B(_471_), .Y(_474_) );
OAI21X1 OAI21X1_237 ( .A(_359_), .B(_471_), .C(_474_), .Y(_1443__2_) );
NAND2X1 NAND2X1_170 ( .A(AXYS_0__3_), .B(_471_), .Y(_475_) );
OAI21X1 OAI21X1_238 ( .A(_366_), .B(_471_), .C(_475_), .Y(_1443__3_) );
NAND2X1 NAND2X1_171 ( .A(AXYS_0__4_), .B(new_wire_71), .Y(_476_) );
OAI21X1 OAI21X1_239 ( .A(_369_), .B(new_wire_71), .C(_476_), .Y(_1443__4_) );
NAND2X1 NAND2X1_172 ( .A(AXYS_0__5_), .B(new_wire_71), .Y(_477_) );
OAI21X1 OAI21X1_240 ( .A(_378_), .B(new_wire_71), .C(_477_), .Y(_1443__5_) );
NAND2X1 NAND2X1_173 ( .A(AXYS_0__6_), .B(new_wire_71), .Y(_478_) );
OAI21X1 OAI21X1_241 ( .A(_383_), .B(new_wire_71), .C(_478_), .Y(_1443__6_) );
NAND2X1 NAND2X1_174 ( .A(AXYS_0__7_), .B(new_wire_71), .Y(_479_) );
OAI21X1 OAI21X1_242 ( .A(_390_), .B(new_wire_71), .C(_479_), .Y(_1443__7_) );
NAND2X1 NAND2X1_175 ( .A(_1094_), .B(_415_), .Y(_480_) );
OAI21X1 OAI21X1_243 ( .A(_1017__bF_buf1), .B(_822__bF_buf4), .C(load_only), .Y(_481_) );
OAI21X1 OAI21X1_244 ( .A(_1101__bF_buf0), .B(_480_), .C(_481_), .Y(_26_) );
NAND3X1 NAND3X1_141 ( .A(_1141_), .B(_1388_), .C(_482_), .Y(_483_) );
OAI21X1 OAI21X1_245 ( .A(_1212_), .B(_1070__bF_buf3), .C(_483_), .Y(_40_) );
NOR2X1 NOR2X1_175 ( .A(new_wire_53), .B(new_wire_54), .Y(_484_) );
OAI21X1 OAI21X1_246 ( .A(_419_), .B(_425_), .C(_484_), .Y(_485_) );
OAI22X1 OAI22X1_40 ( .A(_279_), .B(_1070__bF_buf2), .C(_399_), .D(_485_), .Y(_39_) );
NOR2X1 NOR2X1_176 ( .A(_1358_), .B(_482_), .Y(_486_) );
NAND3X1 NAND3X1_142 ( .A(_1080_), .B(_1331_), .C(_486_), .Y(_487_) );
MUX2X1 MUX2X1_21 ( .A(_1184_), .B(index_y), .S(_1070__bF_buf4), .Y(_488_) );
NAND3X1 NAND3X1_143 ( .A(_1322_), .B(_488_), .C(_487_), .Y(_25_) );
NAND3X1 NAND3X1_144 ( .A(_415_), .B(_426_), .C(_1086_), .Y(_490_) );
NOR2X1 NOR2X1_177 ( .A(_401_), .B(_482_), .Y(_491_) );
OAI21X1 OAI21X1_247 ( .A(_1087_), .B(_492_), .C(_490_), .Y(_493_) );
OAI21X1 OAI21X1_248 ( .A(_825__bF_buf0), .B(_1093_), .C(new_wire_58), .Y(_494_) );
OAI21X1 OAI21X1_249 ( .A(_494_), .B(_495_), .C(_428_), .Y(_496_) );
NOR2X1 NOR2X1_178 ( .A(_496_), .B(_493_), .Y(_497_) );
OAI21X1 OAI21X1_250 ( .A(_1389_), .B(_416_), .C(_497_), .Y(_498_) );
NAND2X1 NAND2X1_176 ( .A(_1070__bF_buf2), .B(_498_), .Y(_499_) );
OAI21X1 OAI21X1_251 ( .A(_489_), .B(_1070__bF_buf2), .C(_499_), .Y(_38__0_) );
NAND2X1 NAND2X1_177 ( .A(_408_), .B(_1095_), .Y(_500_) );
OAI21X1 OAI21X1_252 ( .A(_500_), .B(_1389_), .C(_1070__bF_buf1), .Y(_501_) );
NOR2X1 NOR2X1_179 ( .A(new_wire_54), .B(_1077_), .Y(_502_) );
OAI21X1 OAI21X1_253 ( .A(_426_), .B(_502_), .C(_486_), .Y(_503_) );
OAI21X1 OAI21X1_254 ( .A(_1268_), .B(_495_), .C(_503_), .Y(_504_) );
NOR2X1 NOR2X1_180 ( .A(_501_), .B(_504_), .Y(_505_) );
AOI22X1 AOI22X1_39 ( .A(_128_), .B(_1101__bF_buf1), .C(_505_), .D(_497_), .Y(_38__1_) );
OAI21X1 OAI21X1_255 ( .A(new_wire_58), .B(_1080_), .C(_1086_), .Y(_507_) );
OAI21X1 OAI21X1_256 ( .A(_480_), .B(_507_), .C(_428_), .Y(_508_) );
OAI21X1 OAI21X1_257 ( .A(_1389_), .B(_492_), .C(_397_), .Y(_509_) );
OAI21X1 OAI21X1_258 ( .A(_508_), .B(_509_), .C(_1070__bF_buf0), .Y(_510_) );
OAI21X1 OAI21X1_259 ( .A(_506_), .B(_1070__bF_buf2), .C(_510_), .Y(_23__0_) );
AOI21X1 AOI21X1_79 ( .A(new_wire_54), .B(_486_), .C(_501_), .Y(_511_) );
OAI21X1 OAI21X1_260 ( .A(_1268_), .B(_409_), .C(_511_), .Y(_512_) );
NOR2X1 NOR2X1_181 ( .A(_508_), .B(_512_), .Y(_513_) );
AOI21X1 AOI21X1_80 ( .A(_141_), .B(_1101__bF_buf1), .C(_513_), .Y(_23__1_) );
OAI21X1 OAI21X1_261 ( .A(_1389_), .B(_416_), .C(_433_), .Y(_514_) );
NOR2X1 NOR2X1_182 ( .A(_418_), .B(_416_), .Y(_515_) );
NOR2X1 NOR2X1_183 ( .A(_1080_), .B(_1085_), .Y(_516_) );
NAND3X1 NAND3X1_145 ( .A(_516_), .B(_415_), .C(_502_), .Y(_517_) );
OAI21X1 OAI21X1_262 ( .A(_1274_), .B(_1389_), .C(_517_), .Y(_518_) );
NOR2X1 NOR2X1_184 ( .A(_515_), .B(_518_), .Y(_519_) );
OAI21X1 OAI21X1_263 ( .A(_1188_), .B(_1292_), .C(_519_), .Y(_520_) );
OAI22X1 OAI22X1_41 ( .A(_1183_), .B(_484_), .C(new_wire_56), .D(_1087_), .Y(_521_) );
OR2X2 OR2X2_20 ( .A(_520_), .B(_521_), .Y(_522_) );
OAI21X1 OAI21X1_264 ( .A(_514_), .B(_522_), .C(_1070__bF_buf1), .Y(_523_) );
OAI21X1 OAI21X1_265 ( .A(_338_), .B(_1070__bF_buf3), .C(_523_), .Y(_27_) );
OAI21X1 OAI21X1_266 ( .A(_1072_), .B(_1251_), .C(RDY_bF_buf0), .Y(_524_) );
OR2X2 OR2X2_21 ( .A(_524_), .B(reset), .Y(_525_) );
OAI21X1 OAI21X1_267 ( .A(reset), .B(_524_), .C(IRHOLD_0_), .Y(_526_) );
OAI21X1 OAI21X1_268 ( .A(_104_), .B(_525_), .C(_526_), .Y(_4__0_) );
OAI21X1 OAI21X1_269 ( .A(reset), .B(_524_), .C(IRHOLD_1_), .Y(_527_) );
OAI21X1 OAI21X1_270 ( .A(_118_), .B(_525_), .C(_527_), .Y(_4__1_) );
OAI21X1 OAI21X1_271 ( .A(reset), .B(_524_), .C(IRHOLD_2_), .Y(_528_) );
OAI21X1 OAI21X1_272 ( .A(_978_), .B(_525_), .C(_528_), .Y(_4__2_) );
OAI21X1 OAI21X1_273 ( .A(reset), .B(_524_), .C(IRHOLD_3_), .Y(_529_) );
OAI21X1 OAI21X1_274 ( .A(_1179_), .B(_525_), .C(_529_), .Y(_4__3_) );
MUX2X1 MUX2X1_22 ( .A(_530_), .B(_1019_), .S(_525_), .Y(_4__4_) );
MUX2X1 MUX2X1_23 ( .A(_531_), .B(_119_), .S(_525_), .Y(_4__5_) );
MUX2X1 MUX2X1_24 ( .A(_532_), .B(_1052_), .S(_525_), .Y(_4__6_) );
MUX2X1 MUX2X1_25 ( .A(_533_), .B(_1064_), .S(_525_), .Y(_4__7_) );
OAI21X1 OAI21X1_275 ( .A(_1017__bF_buf3), .B(_822__bF_buf1), .C(new_wire_52), .Y(_534_) );
OAI21X1 OAI21X1_276 ( .A(reset), .B(_534_), .C(new_wire_72), .Y(_5_) );
AOI21X1 AOI21X1_81 ( .A(_1306_), .B(_466_), .C(plp), .Y(_535_) );
OAI21X1 OAI21X1_277 ( .A(_466_), .B(AV), .C(_535_), .Y(_536_) );
NOR2X1 NOR2X1_185 ( .A(clv), .B(_536_), .Y(_537_) );
AOI21X1 AOI21X1_82 ( .A(ADD_6_), .B(plp), .C(_537_), .Y(_538_) );
NOR2X1 NOR2X1_186 ( .A(_539_), .B(_1205_), .Y(_540_) );
NAND2X1 NAND2X1_178 ( .A(DIMUX_6_), .B(_540_), .Y(_541_) );
OAI21X1 OAI21X1_278 ( .A(_1306_), .B(_540_), .C(_541_), .Y(_542_) );
NOR2X1 NOR2X1_187 ( .A(_859__bF_buf2), .B(_1155_), .Y(_543_) );
AOI22X1 AOI22X1_40 ( .A(DIMUX_6_), .B(_1155_), .C(_543_), .D(_542_), .Y(_544_) );
OAI21X1 OAI21X1_279 ( .A(_822__bF_buf3), .B(_538_), .C(_544_), .Y(_10_) );
NAND2X1 NAND2X1_179 ( .A(DIMUX_3_), .B(_1155_), .Y(_545_) );
NOR2X1 NOR2X1_188 ( .A(plp), .B(cld), .Y(_546_) );
OAI21X1 OAI21X1_280 ( .A(D), .B(sed), .C(_546_), .Y(_547_) );
OAI21X1 OAI21X1_281 ( .A(_363_), .B(_324_), .C(_547_), .Y(_548_) );
MUX2X1 MUX2X1_26 ( .A(D), .B(_548_), .S(_822__bF_buf3), .Y(_549_) );
OAI21X1 OAI21X1_282 ( .A(_1155_), .B(_549_), .C(_545_), .Y(_3_) );
NAND2X1 NAND2X1_180 ( .A(new_wire_61), .B(_470_), .Y(_550_) );
NAND2X1 NAND2X1_181 ( .A(AXYS_2__0_), .B(_550_), .Y(_551_) );
OAI21X1 OAI21X1_283 ( .A(_345_), .B(_550_), .C(_551_), .Y(_1444__0_) );
NAND2X1 NAND2X1_182 ( .A(AXYS_2__1_), .B(_550_), .Y(_552_) );
OAI21X1 OAI21X1_284 ( .A(_354_), .B(_550_), .C(_552_), .Y(_1444__1_) );
NAND2X1 NAND2X1_183 ( .A(AXYS_2__2_), .B(_550_), .Y(_553_) );
OAI21X1 OAI21X1_285 ( .A(_359_), .B(_550_), .C(_553_), .Y(_1444__2_) );
NAND2X1 NAND2X1_184 ( .A(AXYS_2__3_), .B(_550_), .Y(_554_) );
OAI21X1 OAI21X1_286 ( .A(_366_), .B(_550_), .C(_554_), .Y(_1444__3_) );
NAND2X1 NAND2X1_185 ( .A(AXYS_2__4_), .B(new_wire_73), .Y(_555_) );
OAI21X1 OAI21X1_287 ( .A(_369_), .B(new_wire_73), .C(_555_), .Y(_1444__4_) );
NAND2X1 NAND2X1_186 ( .A(AXYS_2__5_), .B(new_wire_73), .Y(_556_) );
OAI21X1 OAI21X1_288 ( .A(_378_), .B(new_wire_73), .C(_556_), .Y(_1444__5_) );
NAND2X1 NAND2X1_187 ( .A(AXYS_2__6_), .B(new_wire_73), .Y(_557_) );
OAI21X1 OAI21X1_289 ( .A(_383_), .B(new_wire_73), .C(_557_), .Y(_1444__6_) );
NAND2X1 NAND2X1_188 ( .A(AXYS_2__7_), .B(new_wire_73), .Y(_558_) );
OAI21X1 OAI21X1_290 ( .A(_390_), .B(new_wire_73), .C(_558_), .Y(_1444__7_) );
OAI21X1 OAI21X1_291 ( .A(new_wire_61), .B(_155__bF_buf0), .C(load_reg), .Y(_560_) );
AOI21X1 AOI21X1_83 ( .A(_560_), .B(_86_), .C(_559_), .Y(_561_) );
NAND2X1 NAND2X1_189 ( .A(_86_), .B(_560_), .Y(_562_) );
OAI21X1 OAI21X1_292 ( .A(_318_), .B(_562_), .C(_324_), .Y(_563_) );
AOI21X1 AOI21X1_84 ( .A(_387_), .B(plp), .C(_822__bF_buf3), .Y(_564_) );
OAI21X1 OAI21X1_293 ( .A(_561_), .B(_563_), .C(_564_), .Y(_565_) );
OAI21X1 OAI21X1_294 ( .A(_539_), .B(_1205_), .C(_330_), .Y(_566_) );
NAND2X1 NAND2X1_190 ( .A(N), .B(_543_), .Y(_567_) );
OAI21X1 OAI21X1_295 ( .A(_540_), .B(_567_), .C(_1192_), .Y(_568_) );
AOI21X1 AOI21X1_85 ( .A(DIMUX_7_), .B(_566_), .C(_568_), .Y(_569_) );
AOI22X1 AOI22X1_41 ( .A(_559_), .B(_283_), .C(_569_), .D(_565_), .Y(_8_) );
NAND3X1 NAND3X1_146 ( .A(_86_), .B(_539_), .C(_560_), .Y(_571_) );
AND2X2 AND2X2_44 ( .A(_571_), .B(AZ), .Y(_572_) );
OAI21X1 OAI21X1_296 ( .A(_1303_), .B(_571_), .C(_324_), .Y(_573_) );
AOI21X1 AOI21X1_86 ( .A(_931_), .B(plp), .C(_822__bF_buf3), .Y(_574_) );
OAI21X1 OAI21X1_297 ( .A(_572_), .B(_573_), .C(_574_), .Y(_575_) );
OAI21X1 OAI21X1_298 ( .A(_118_), .B(_330_), .C(_1192_), .Y(_576_) );
AOI21X1 AOI21X1_87 ( .A(_543_), .B(Z), .C(_576_), .Y(_577_) );
AOI22X1 AOI22X1_42 ( .A(_570_), .B(_283_), .C(_577_), .D(_575_), .Y(_11_) );
NOR2X1 NOR2X1_189 ( .A(_87_), .B(_1192_), .Y(_578_) );
NAND3X1 NAND3X1_147 ( .A(_86_), .B(_87_), .C(_466_), .Y(_579_) );
NOR2X1 NOR2X1_190 ( .A(plp), .B(clc), .Y(_580_) );
OAI21X1 OAI21X1_299 ( .A(C), .B(sec), .C(_580_), .Y(_581_) );
OAI21X1 OAI21X1_300 ( .A(_904_), .B(_324_), .C(_581_), .Y(_582_) );
NOR2X1 NOR2X1_191 ( .A(write_back), .B(_822__bF_buf3), .Y(_583_) );
OAI21X1 OAI21X1_301 ( .A(_579_), .B(_582_), .C(_583_), .Y(_584_) );
AOI21X1 AOI21X1_88 ( .A(_370_), .B(_579_), .C(_584_), .Y(_585_) );
OAI21X1 OAI21X1_302 ( .A(_79_), .B(_583_), .C(_330_), .Y(_586_) );
OAI22X1 OAI22X1_42 ( .A(DIMUX_0_), .B(_330_), .C(_586_), .D(_585_), .Y(_587_) );
NAND2X1 NAND2X1_191 ( .A(CO), .B(_578_), .Y(_588_) );
OAI21X1 OAI21X1_303 ( .A(_578_), .B(_587_), .C(_588_), .Y(_2_) );
NOR2X1 NOR2X1_192 ( .A(new_wire_62), .B(_342_), .Y(_589_) );
MUX2X1 MUX2X1_27 ( .A(_345_), .B(_158_), .S(_589_), .Y(_1445__0_) );
MUX2X1 MUX2X1_28 ( .A(_354_), .B(_181_), .S(_589_), .Y(_1445__1_) );
MUX2X1 MUX2X1_29 ( .A(_359_), .B(_194_), .S(_589_), .Y(_1445__2_) );
MUX2X1 MUX2X1_30 ( .A(_366_), .B(_207_), .S(_589_), .Y(_1445__3_) );
MUX2X1 MUX2X1_31 ( .A(_369_), .B(_220_), .S(_589_), .Y(_1445__4_) );
MUX2X1 MUX2X1_32 ( .A(_378_), .B(_234_), .S(_589_), .Y(_1445__5_) );
MUX2X1 MUX2X1_33 ( .A(_383_), .B(_247_), .S(_589_), .Y(_1445__6_) );
MUX2X1 MUX2X1_34 ( .A(_390_), .B(_260_), .S(_589_), .Y(_1445__7_) );
NAND2X1 NAND2X1_192 ( .A(new_wire_9), .B(DI[7]), .Y(_590_) );
OAI21X1 OAI21X1_304 ( .A(new_wire_9), .B(_275_), .C(_590_), .Y(_15_) );
NOR2X1 NOR2X1_193 ( .A(_95_), .B(_270_), .Y(_591_) );
AOI21X1 AOI21X1_89 ( .A(_157_), .B(_162_), .C(_591_), .Y(_592_) );
NOR2X1 NOR2X1_194 ( .A(_337_), .B(_94_), .Y(_593_) );
NAND3X1 NAND3X1_148 ( .A(_330_), .B(_136_), .C(_593_), .Y(_594_) );
NOR2X1 NOR2X1_195 ( .A(_121_), .B(_594_), .Y(_595_) );
OAI21X1 OAI21X1_305 ( .A(_809__bF_buf2), .B(_1071_), .C(_1211_), .Y(_596_) );
OR2X2 OR2X2_22 ( .A(_596_), .B(_91_), .Y(_597_) );
NOR2X1 NOR2X1_196 ( .A(_796_), .B(_911_), .Y(_598_) );
OAI21X1 OAI21X1_306 ( .A(_795__bF_buf3), .B(_1071_), .C(_598_), .Y(_599_) );
NOR2X1 NOR2X1_197 ( .A(_597_), .B(_599_), .Y(_600_) );
OAI21X1 OAI21X1_307 ( .A(_809__bF_buf2), .B(_1138_), .C(_1109_), .Y(_601_) );
OAI21X1 OAI21X1_308 ( .A(_795__bF_buf0), .B(_1236_), .C(_1115_), .Y(_602_) );
NOR2X1 NOR2X1_198 ( .A(_602_), .B(_601_), .Y(_603_) );
NAND3X1 NAND3X1_149 ( .A(_603_), .B(_600_), .C(_595_), .Y(_604_) );
OAI21X1 OAI21X1_309 ( .A(_799__bF_buf4), .B(new_wire_57), .C(_80_), .Y(_605_) );
OR2X2 OR2X2_23 ( .A(_605_), .B(_849__bF_buf2), .Y(_606_) );
NAND2X1 NAND2X1_193 ( .A(new_wire_31), .B(_920_), .Y(_607_) );
NAND3X1 NAND3X1_150 ( .A(_847_), .B(_607_), .C(_1197_), .Y(_608_) );
OAI21X1 OAI21X1_310 ( .A(_799__bF_buf4), .B(_1138_), .C(_1320_), .Y(_609_) );
NOR2X1 NOR2X1_199 ( .A(_608_), .B(_609_), .Y(_610_) );
NAND2X1 NAND2X1_194 ( .A(_610_), .B(_591_), .Y(_611_) );
OR2X2 OR2X2_24 ( .A(_611_), .B(_606_), .Y(_612_) );
OR2X2 OR2X2_25 ( .A(_612_), .B(_604_), .Y(_613_) );
AOI22X1 AOI22X1_43 ( .A(ADD_0_), .B(_849__bF_buf1), .C(DIMUX_0_), .D(_609_), .Y(_615_) );
NOR2X1 NOR2X1_200 ( .A(_608_), .B(_605_), .Y(_616_) );
OAI21X1 OAI21X1_311 ( .A(_614_), .B(_616_), .C(_615_), .Y(_617_) );
AOI21X1 AOI21X1_90 ( .A(_604_), .B(ADD_0_), .C(_617_), .Y(_618_) );
OAI21X1 OAI21X1_312 ( .A(_905_), .B(_613_), .C(_618_), .Y(_619_) );
OR2X2 OR2X2_26 ( .A(_619_), .B(_592_), .Y(_1439__0_) );
OAI21X1 OAI21X1_313 ( .A(_920_), .B(_1196_), .C(new_wire_31), .Y(_620_) );
NAND2X1 NAND2X1_195 ( .A(_621_), .B(_543_), .Y(_622_) );
AOI21X1 AOI21X1_91 ( .A(new_wire_31), .B(_838_), .C(_1312_), .Y(_623_) );
NAND3X1 NAND3X1_151 ( .A(_166_), .B(_623_), .C(_598_), .Y(_624_) );
NOR2X1 NOR2X1_201 ( .A(_622_), .B(_624_), .Y(_625_) );
OR2X2 OR2X2_27 ( .A(_922_), .B(new_wire_46), .Y(_626_) );
NAND2X1 NAND2X1_196 ( .A(_107_), .B(_164_), .Y(_627_) );
OR2X2 OR2X2_28 ( .A(_626_), .B(_627_), .Y(_628_) );
NOR2X1 NOR2X1_202 ( .A(_122_), .B(_628_), .Y(_629_) );
NAND3X1 NAND3X1_152 ( .A(_620_), .B(_625_), .C(_629_), .Y(_630_) );
NOR2X1 NOR2X1_203 ( .A(_807_), .B(_96_), .Y(_631_) );
NAND3X1 NAND3X1_153 ( .A(_136_), .B(_620_), .C(_114_), .Y(_632_) );
NOR2X1 NOR2X1_204 ( .A(_632_), .B(_108_), .Y(_633_) );
NOR2X1 NOR2X1_205 ( .A(_328_), .B(_1072_), .Y(_634_) );
OAI21X1 OAI21X1_314 ( .A(_621_), .B(_634_), .C(_543_), .Y(_635_) );
NOR2X1 NOR2X1_206 ( .A(_1336_), .B(_1099_), .Y(_636_) );
NOR2X1 NOR2X1_207 ( .A(_1416_), .B(new_wire_59), .Y(_637_) );
NAND3X1 NAND3X1_154 ( .A(_110_), .B(_637_), .C(_636_), .Y(_638_) );
NOR2X1 NOR2X1_208 ( .A(_635_), .B(_638_), .Y(_639_) );
NAND3X1 NAND3X1_155 ( .A(_631_), .B(_633_), .C(_639_), .Y(_640_) );
NOR2X1 NOR2X1_209 ( .A(_596_), .B(_601_), .Y(_641_) );
NOR2X1 NOR2X1_210 ( .A(_337_), .B(_609_), .Y(_642_) );
AND2X2 AND2X2_45 ( .A(_642_), .B(_641_), .Y(_643_) );
NAND3X1 NAND3X1_156 ( .A(_1197_), .B(_1115_), .C(_1150_), .Y(_644_) );
NAND3X1 NAND3X1_157 ( .A(_925_), .B(_1114_), .C(_1404_), .Y(_645_) );
NOR2X1 NOR2X1_211 ( .A(_644_), .B(_645_), .Y(_646_) );
NOR2X1 NOR2X1_212 ( .A(_605_), .B(_647_), .Y(_648_) );
NAND3X1 NAND3X1_158 ( .A(_646_), .B(_648_), .C(_643_), .Y(_649_) );
AOI21X1 AOI21X1_92 ( .A(_630_), .B(_640_), .C(_649_), .Y(_650_) );
NOR2X1 NOR2X1_213 ( .A(_1017__bF_buf2), .B(_650_), .Y(_651_) );
OAI21X1 OAI21X1_315 ( .A(_619_), .B(_592_), .C(_651__bF_buf2), .Y(_652_) );
OAI21X1 OAI21X1_316 ( .A(_614_), .B(_651__bF_buf2), .C(_652_), .Y(_1__0_) );
AOI21X1 AOI21X1_93 ( .A(_180_), .B(_185_), .C(_591_), .Y(_653_) );
AOI22X1 AOI22X1_44 ( .A(ADD_1_), .B(_849__bF_buf1), .C(DIMUX_1_), .D(_609_), .Y(_655_) );
OAI21X1 OAI21X1_317 ( .A(_654_), .B(_616_), .C(_655_), .Y(_656_) );
AOI21X1 AOI21X1_94 ( .A(_604_), .B(ADD_1_), .C(_656_), .Y(_657_) );
OAI21X1 OAI21X1_318 ( .A(_933_), .B(_613_), .C(_657_), .Y(_658_) );
OR2X2 OR2X2_29 ( .A(_658_), .B(_653_), .Y(_1439__1_) );
OAI21X1 OAI21X1_319 ( .A(_658_), .B(_653_), .C(_651__bF_buf4), .Y(_659_) );
OAI21X1 OAI21X1_320 ( .A(_654_), .B(_651__bF_buf4), .C(_659_), .Y(_1__1_) );
AOI21X1 AOI21X1_95 ( .A(_193_), .B(_198_), .C(_591_), .Y(_660_) );
AOI22X1 AOI22X1_45 ( .A(new_wire_51), .B(_849__bF_buf3), .C(DIMUX_2_), .D(_609_), .Y(_661_) );
OAI21X1 OAI21X1_321 ( .A(_958_), .B(_616_), .C(_661_), .Y(_662_) );
AOI21X1 AOI21X1_96 ( .A(_604_), .B(new_wire_51), .C(_662_), .Y(_663_) );
OAI21X1 OAI21X1_322 ( .A(_956_), .B(_613_), .C(_663_), .Y(_664_) );
OR2X2 OR2X2_30 ( .A(_664_), .B(_660_), .Y(_1439__2_) );
OAI21X1 OAI21X1_323 ( .A(_664_), .B(_660_), .C(_651__bF_buf0), .Y(_665_) );
OAI21X1 OAI21X1_324 ( .A(_958_), .B(_651__bF_buf0), .C(_665_), .Y(_1__2_) );
AOI21X1 AOI21X1_97 ( .A(_206_), .B(_211_), .C(_591_), .Y(_666_) );
AOI22X1 AOI22X1_46 ( .A(ADD_3_), .B(_849__bF_buf3), .C(DIMUX_3_), .D(_609_), .Y(_667_) );
OAI21X1 OAI21X1_325 ( .A(_946_), .B(_616_), .C(_667_), .Y(_668_) );
AOI21X1 AOI21X1_98 ( .A(_604_), .B(new_wire_50), .C(_668_), .Y(_669_) );
OAI21X1 OAI21X1_326 ( .A(_944_), .B(_613_), .C(_669_), .Y(_670_) );
OR2X2 OR2X2_31 ( .A(_670_), .B(_666_), .Y(_1439__3_) );
OAI21X1 OAI21X1_327 ( .A(_670_), .B(_666_), .C(_651__bF_buf0), .Y(_671_) );
OAI21X1 OAI21X1_328 ( .A(_946_), .B(_651__bF_buf0), .C(_671_), .Y(_1__3_) );
AOI21X1 AOI21X1_99 ( .A(_219_), .B(_224_), .C(_591_), .Y(_672_) );
AOI22X1 AOI22X1_47 ( .A(ADD_4_), .B(_849__bF_buf1), .C(DIMUX_4_), .D(_609_), .Y(_673_) );
OAI21X1 OAI21X1_329 ( .A(_874_), .B(_616_), .C(_673_), .Y(_674_) );
AOI21X1 AOI21X1_100 ( .A(_604_), .B(ADD_4_), .C(_674_), .Y(_675_) );
OAI21X1 OAI21X1_330 ( .A(_872_), .B(_613_), .C(_675_), .Y(_676_) );
OR2X2 OR2X2_32 ( .A(_676_), .B(_672_), .Y(_1439__4_) );
OAI21X1 OAI21X1_331 ( .A(_676_), .B(_672_), .C(_651__bF_buf1), .Y(_677_) );
OAI21X1 OAI21X1_332 ( .A(_874_), .B(_651__bF_buf1), .C(_677_), .Y(_1__4_) );
AOI21X1 AOI21X1_101 ( .A(_233_), .B(_238_), .C(_591_), .Y(_678_) );
AOI22X1 AOI22X1_48 ( .A(ADD_5_), .B(_849__bF_buf1), .C(DIMUX_5_), .D(_609_), .Y(_679_) );
OAI21X1 OAI21X1_333 ( .A(_862_), .B(_616_), .C(_679_), .Y(_680_) );
AOI21X1 AOI21X1_102 ( .A(_604_), .B(ADD_5_), .C(_680_), .Y(_681_) );
OAI21X1 OAI21X1_334 ( .A(_860_), .B(_613_), .C(_681_), .Y(_682_) );
OR2X2 OR2X2_33 ( .A(_682_), .B(_678_), .Y(_1439__5_) );
OAI21X1 OAI21X1_335 ( .A(_682_), .B(_678_), .C(_651__bF_buf1), .Y(_683_) );
OAI21X1 OAI21X1_336 ( .A(_862_), .B(_651__bF_buf2), .C(_683_), .Y(_1__5_) );
AOI21X1 AOI21X1_103 ( .A(_246_), .B(_251_), .C(_591_), .Y(_684_) );
AOI22X1 AOI22X1_49 ( .A(new_wire_48), .B(_849__bF_buf2), .C(DIMUX_6_), .D(new_wire_76), .Y(_685_) );
OAI21X1 OAI21X1_337 ( .A(_895_), .B(_616_), .C(_685_), .Y(_686_) );
AOI21X1 AOI21X1_104 ( .A(_604_), .B(new_wire_48), .C(_686_), .Y(_687_) );
OAI21X1 OAI21X1_338 ( .A(_893_), .B(_613_), .C(_687_), .Y(_688_) );
OR2X2 OR2X2_34 ( .A(_688_), .B(_684_), .Y(_1439__6_) );
OAI21X1 OAI21X1_339 ( .A(_688_), .B(_684_), .C(_651__bF_buf0), .Y(_689_) );
OAI21X1 OAI21X1_340 ( .A(_895_), .B(_651__bF_buf0), .C(_689_), .Y(_1__6_) );
AOI21X1 AOI21X1_105 ( .A(_259_), .B(_264_), .C(new_wire_74), .Y(_690_) );
AOI22X1 AOI22X1_50 ( .A(ADD_7_), .B(_849__bF_buf2), .C(DIMUX_7_), .D(new_wire_76), .Y(_691_) );
OAI21X1 OAI21X1_341 ( .A(_885_), .B(_616_), .C(_691_), .Y(_692_) );
AOI21X1 AOI21X1_106 ( .A(new_wire_75), .B(ADD_7_), .C(_692_), .Y(_693_) );
OAI21X1 OAI21X1_342 ( .A(_883_), .B(_613_), .C(_693_), .Y(_694_) );
OR2X2 OR2X2_35 ( .A(_694_), .B(_690_), .Y(_1439__7_) );
OAI21X1 OAI21X1_343 ( .A(_694_), .B(_690_), .C(_651__bF_buf1), .Y(_695_) );
OAI21X1 OAI21X1_344 ( .A(_885_), .B(_651__bF_buf2), .C(_695_), .Y(_1__7_) );
OAI21X1 OAI21X1_345 ( .A(_88_), .B(_283_), .C(ABH_0_), .Y(_696_) );
AOI21X1 AOI21X1_107 ( .A(_608_), .B(new_wire_49), .C(_120_), .Y(_697_) );
NAND3X1 NAND3X1_159 ( .A(_696_), .B(_697_), .C(new_wire_74), .Y(_698_) );
OAI21X1 OAI21X1_346 ( .A(_104_), .B(_600_), .C(_595_), .Y(_699_) );
NOR2X1 NOR2X1_214 ( .A(_698_), .B(_699_), .Y(_700_) );
OAI21X1 OAI21X1_347 ( .A(_1008_), .B(new_wire_77), .C(_700_), .Y(_1439__8_) );
NAND2X1 NAND2X1_197 ( .A(_1439__8_), .B(_651__bF_buf4), .Y(_701_) );
OAI21X1 OAI21X1_348 ( .A(_1006_), .B(_651__bF_buf4), .C(_701_), .Y(_0__0_) );
OAI21X1 OAI21X1_349 ( .A(_849__bF_buf3), .B(_605_), .C(ABH_1_), .Y(_704_) );
OAI21X1 OAI21X1_350 ( .A(_931_), .B(_703_), .C(_704_), .Y(_705_) );
AOI21X1 AOI21X1_108 ( .A(_702_), .B(DIMUX_1_), .C(_705_), .Y(_706_) );
OAI21X1 OAI21X1_351 ( .A(_996_), .B(new_wire_77), .C(_706_), .Y(_1439__9_) );
NAND2X1 NAND2X1_198 ( .A(_1439__9_), .B(_651__bF_buf2), .Y(_707_) );
OAI21X1 OAI21X1_352 ( .A(_994_), .B(_651__bF_buf2), .C(_707_), .Y(_0__1_) );
OAI21X1 OAI21X1_353 ( .A(_849__bF_buf3), .B(_605_), .C(ABH_2_), .Y(_708_) );
OAI21X1 OAI21X1_354 ( .A(_360_), .B(_703_), .C(_708_), .Y(_709_) );
AOI21X1 AOI21X1_109 ( .A(_702_), .B(DIMUX_2_), .C(_709_), .Y(_710_) );
OAI21X1 OAI21X1_355 ( .A(_983_), .B(new_wire_77), .C(_710_), .Y(_1439__10_) );
NAND2X1 NAND2X1_199 ( .A(_1439__10_), .B(_651__bF_buf1), .Y(_711_) );
OAI21X1 OAI21X1_356 ( .A(_981_), .B(_651__bF_buf1), .C(_711_), .Y(_0__2_) );
OAI21X1 OAI21X1_357 ( .A(_849__bF_buf3), .B(_605_), .C(ABH_3_), .Y(_712_) );
OAI21X1 OAI21X1_358 ( .A(_363_), .B(_703_), .C(_712_), .Y(_713_) );
AOI21X1 AOI21X1_110 ( .A(_702_), .B(DIMUX_3_), .C(_713_), .Y(_714_) );
OAI21X1 OAI21X1_359 ( .A(_972_), .B(new_wire_77), .C(_714_), .Y(_1439__11_) );
NAND2X1 NAND2X1_200 ( .A(_1439__11_), .B(_651__bF_buf4), .Y(_715_) );
OAI21X1 OAI21X1_360 ( .A(_970_), .B(_651__bF_buf4), .C(_715_), .Y(_0__3_) );
OAI22X1 OAI22X1_43 ( .A(_367_), .B(_703_), .C(_1019_), .D(_600_), .Y(_716_) );
AOI21X1 AOI21X1_111 ( .A(ABH_4_), .B(_606_), .C(_716_), .Y(_717_) );
OAI21X1 OAI21X1_361 ( .A(_1016_), .B(new_wire_77), .C(_717_), .Y(_1439__12_) );
NAND2X1 NAND2X1_201 ( .A(_1439__12_), .B(_651__bF_buf4), .Y(_718_) );
OAI21X1 OAI21X1_362 ( .A(_1020_), .B(_651__bF_buf3), .C(_718_), .Y(_0__4_) );
OAI21X1 OAI21X1_363 ( .A(_849__bF_buf2), .B(_605_), .C(ABH_5_), .Y(_719_) );
OAI21X1 OAI21X1_364 ( .A(_846_), .B(_703_), .C(_719_), .Y(_720_) );
AOI21X1 AOI21X1_112 ( .A(_702_), .B(DIMUX_5_), .C(_720_), .Y(_721_) );
OAI21X1 OAI21X1_365 ( .A(_787_), .B(new_wire_77), .C(_721_), .Y(_1439__13_) );
NAND2X1 NAND2X1_202 ( .A(_1439__13_), .B(_651__bF_buf3), .Y(_722_) );
OAI21X1 OAI21X1_366 ( .A(_226_), .B(_651__bF_buf3), .C(_722_), .Y(_0__5_) );
OAI21X1 OAI21X1_367 ( .A(_849__bF_buf4), .B(_605_), .C(ABH_6_), .Y(_724_) );
OAI21X1 OAI21X1_368 ( .A(_384_), .B(_703_), .C(_724_), .Y(_725_) );
AOI21X1 AOI21X1_113 ( .A(_702_), .B(DIMUX_6_), .C(_725_), .Y(_726_) );
OAI21X1 OAI21X1_369 ( .A(_723_), .B(new_wire_77), .C(_726_), .Y(_1439__14_) );
NAND2X1 NAND2X1_203 ( .A(_1439__14_), .B(_651__bF_buf3), .Y(_727_) );
OAI21X1 OAI21X1_370 ( .A(_1049_), .B(_651__bF_buf3), .C(_727_), .Y(_0__6_) );
OAI22X1 OAI22X1_44 ( .A(_387_), .B(_703_), .C(_1064_), .D(_600_), .Y(_728_) );
AOI21X1 AOI21X1_114 ( .A(ABH_7_), .B(_606_), .C(_728_), .Y(_729_) );
OAI21X1 OAI21X1_371 ( .A(_1059_), .B(new_wire_77), .C(_729_), .Y(_1439__15_) );
NAND2X1 NAND2X1_204 ( .A(_1439__15_), .B(_651__bF_buf3), .Y(_730_) );
OAI21X1 OAI21X1_372 ( .A(_1061_), .B(_651__bF_buf3), .C(_730_), .Y(_0__7_) );
OAI21X1 OAI21X1_373 ( .A(_905_), .B(_820_), .C(_910_), .Y(_731_) );
NAND2X1 NAND2X1_205 ( .A(_918_), .B(_927_), .Y(_732_) );
NOR2X1 NOR2X1_215 ( .A(_732_), .B(_731_), .Y(_733_) );
OAI21X1 OAI21X1_374 ( .A(_904_), .B(new_wire_33), .C(_909_), .Y(_735_) );
OAI21X1 OAI21X1_375 ( .A(_735_), .B(_734_), .C(_732_), .Y(_736_) );
NAND2X1 NAND2X1_206 ( .A(RDY_bF_buf7), .B(_736_), .Y(_737_) );
OAI22X1 OAI22X1_45 ( .A(new_wire_2), .B(_905_), .C(_733_), .D(_737_), .Y(_9__0_) );
NOR2X1 NOR2X1_216 ( .A(_940_), .B(_928_), .Y(_738_) );
NAND2X1 NAND2X1_207 ( .A(RDY_bF_buf3), .B(_1031_), .Y(_739_) );
OAI22X1 OAI22X1_46 ( .A(RDY_bF_buf3), .B(_933_), .C(_738_), .D(_739_), .Y(_9__1_) );
OAI21X1 OAI21X1_376 ( .A(_956_), .B(_820_), .C(_962_), .Y(_741_) );
NOR2X1 NOR2X1_217 ( .A(_741_), .B(_740_), .Y(_742_) );
NAND3X1 NAND3X1_160 ( .A(_940_), .B(_741_), .C(_928_), .Y(_743_) );
NAND2X1 NAND2X1_208 ( .A(RDY_bF_buf3), .B(_743_), .Y(_744_) );
OAI22X1 OAI22X1_47 ( .A(RDY_bF_buf6), .B(_956_), .C(_744_), .D(_742_), .Y(_9__2_) );
NOR2X1 NOR2X1_218 ( .A(_1035_), .B(_1032_), .Y(_745_) );
AND2X2 AND2X2_46 ( .A(_743_), .B(_745_), .Y(_746_) );
OAI21X1 OAI21X1_377 ( .A(_745_), .B(_743_), .C(RDY_bF_buf3), .Y(_747_) );
OAI22X1 OAI22X1_48 ( .A(RDY_bF_buf3), .B(_944_), .C(_746_), .D(_747_), .Y(_9__3_) );
OAI21X1 OAI21X1_378 ( .A(_872_), .B(_820_), .C(_878_), .Y(_748_) );
NOR2X1 NOR2X1_219 ( .A(_745_), .B(_743_), .Y(_749_) );
AOI21X1 AOI21X1_115 ( .A(_749_), .B(_748_), .C(_1017__bF_buf4), .Y(_750_) );
OAI21X1 OAI21X1_379 ( .A(_748_), .B(_749_), .C(_750_), .Y(_751_) );
OAI21X1 OAI21X1_380 ( .A(RDY_bF_buf6), .B(_872_), .C(_751_), .Y(_9__4_) );
OAI21X1 OAI21X1_381 ( .A(_860_), .B(_820_), .C(_867_), .Y(_752_) );
AOI21X1 AOI21X1_116 ( .A(_749_), .B(_748_), .C(_752_), .Y(_753_) );
NOR3X1 NOR3X1_15 ( .A(_745_), .B(_754_), .C(_743_), .Y(_755_) );
OR2X2 OR2X2_36 ( .A(_755_), .B(_1017__bF_buf4), .Y(_756_) );
OAI22X1 OAI22X1_49 ( .A(RDY_bF_buf3), .B(_860_), .C(_753_), .D(_756_), .Y(_9__5_) );
OAI21X1 OAI21X1_382 ( .A(_893_), .B(_820_), .C(_899_), .Y(_757_) );
AOI21X1 AOI21X1_117 ( .A(_755_), .B(_757_), .C(_1017__bF_buf4), .Y(_758_) );
OAI21X1 OAI21X1_383 ( .A(_757_), .B(_755_), .C(_758_), .Y(_759_) );
OAI21X1 OAI21X1_384 ( .A(new_wire_6), .B(_893_), .C(_759_), .Y(_9__6_) );
OAI21X1 OAI21X1_385 ( .A(_883_), .B(_820_), .C(_889_), .Y(_760_) );
AOI21X1 AOI21X1_118 ( .A(_755_), .B(_757_), .C(_760_), .Y(_761_) );
NAND3X1 NAND3X1_161 ( .A(_760_), .B(_757_), .C(_755_), .Y(_762_) );
NAND2X1 NAND2X1_209 ( .A(new_wire_2), .B(_762_), .Y(_763_) );
OAI22X1 OAI22X1_50 ( .A(new_wire_2), .B(_883_), .C(_761_), .D(_763_), .Y(_9__7_) );
OAI21X1 OAI21X1_386 ( .A(_1008_), .B(new_wire_36), .C(_1012_), .Y(_764_) );
OAI21X1 OAI21X1_387 ( .A(_901_), .B(_964_), .C(_764_), .Y(_765_) );
NAND3X1 NAND3X1_162 ( .A(_963_), .B(_1030_), .C(_740_), .Y(_766_) );
OR2X2 OR2X2_37 ( .A(_766_), .B(_764_), .Y(_767_) );
NAND3X1 NAND3X1_163 ( .A(RDY_bF_buf6), .B(_765_), .C(_767_), .Y(_768_) );
NAND2X1 NAND2X1_210 ( .A(_1017__bF_buf4), .B(_1008_), .Y(_769_) );
AND2X2 AND2X2_47 ( .A(_768_), .B(_769_), .Y(_9__8_) );
OAI21X1 OAI21X1_388 ( .A(_996_), .B(new_wire_36), .C(_1000_), .Y(_770_) );
NOR2X1 NOR2X1_220 ( .A(_901_), .B(_964_), .Y(_771_) );
AOI21X1 AOI21X1_119 ( .A(_771_), .B(_764_), .C(_770_), .Y(_772_) );
OAI21X1 OAI21X1_389 ( .A(_773_), .B(_766_), .C(RDY_bF_buf6), .Y(_774_) );
OAI22X1 OAI22X1_51 ( .A(RDY_bF_buf6), .B(_996_), .C(_772_), .D(_774_), .Y(_9__9_) );
OAI21X1 OAI21X1_390 ( .A(_983_), .B(new_wire_36), .C(_987_), .Y(_775_) );
NOR2X1 NOR2X1_221 ( .A(_773_), .B(_766_), .Y(_776_) );
NOR2X1 NOR2X1_222 ( .A(_775_), .B(_776_), .Y(_777_) );
NAND2X1 NAND2X1_211 ( .A(_1013_), .B(_771_), .Y(_779_) );
OAI21X1 OAI21X1_391 ( .A(_778_), .B(_779_), .C(RDY_bF_buf6), .Y(_780_) );
OAI22X1 OAI22X1_52 ( .A(new_wire_3), .B(_983_), .C(_780_), .D(_777_), .Y(_9__10_) );
OAI21X1 OAI21X1_392 ( .A(_972_), .B(new_wire_36), .C(_976_), .Y(_781_) );
AOI21X1 AOI21X1_120 ( .A(_776_), .B(_775_), .C(_781_), .Y(_782_) );
OAI21X1 OAI21X1_393 ( .A(_1014_), .B(_766_), .C(new_wire_3), .Y(_783_) );
OAI22X1 OAI22X1_53 ( .A(new_wire_3), .B(_972_), .C(_783_), .D(_782_), .Y(_9__11_) );
NOR2X1 NOR2X1_223 ( .A(_1028_), .B(_1015_), .Y(_784_) );
OAI21X1 OAI21X1_394 ( .A(_785_), .B(_1043_), .C(new_wire_6), .Y(_786_) );
OAI22X1 OAI22X1_54 ( .A(new_wire_6), .B(_1016_), .C(_784_), .D(_786_), .Y(_9__12_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf8), .D(_1443__0_), .Q(AXYS_0__0_) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf5), .D(_1443__1_), .Q(AXYS_0__1_) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf11), .D(_1443__2_), .Q(AXYS_0__2_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf7), .D(_1443__3_), .Q(AXYS_0__3_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf5), .D(_1443__4_), .Q(AXYS_0__4_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf8), .D(_1443__5_), .Q(AXYS_0__5_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf8), .D(_1443__6_), .Q(AXYS_0__6_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf11), .D(_1443__7_), .Q(AXYS_0__7_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf5), .D(_1442__0_), .Q(AXYS_1__0_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf7), .D(_1442__1_), .Q(AXYS_1__1_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf11), .D(_1442__2_), .Q(AXYS_1__2_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf8), .D(_1442__3_), .Q(AXYS_1__3_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf5), .D(_1442__4_), .Q(AXYS_1__4_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf8), .D(_1442__5_), .Q(AXYS_1__5_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf8), .D(_1442__6_), .Q(AXYS_1__6_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf11), .D(_1442__7_), .Q(AXYS_1__7_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf8), .D(_1445__0_), .Q(AXYS_3__0_) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf5), .D(_1445__1_), .Q(AXYS_3__1_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf11), .D(_1445__2_), .Q(AXYS_3__2_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf11), .D(_1445__3_), .Q(AXYS_3__3_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf5), .D(_1445__4_), .Q(AXYS_3__4_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf11), .D(_1445__5_), .Q(AXYS_3__5_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf8), .D(_1445__6_), .Q(AXYS_3__6_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf11), .D(_1445__7_), .Q(AXYS_3__7_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(new_wire_13), .D(_1444__0_), .Q(AXYS_2__0_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf5), .D(_1444__1_), .Q(AXYS_2__1_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(new_wire_10), .D(_1444__2_), .Q(AXYS_2__2_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf6), .D(_1444__3_), .Q(AXYS_2__3_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf5), .D(_1444__4_), .Q(AXYS_2__4_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(new_wire_16), .D(_1444__5_), .Q(AXYS_2__5_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(new_wire_13), .D(_1444__6_), .Q(AXYS_2__6_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(new_wire_10), .D(_1444__7_), .Q(AXYS_2__7_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf7), .D(_7_), .Q(NMI_edge) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(new_wire_10), .D(NMI), .Q(NMI_1) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf10), .D(_22__0_), .Q(cond_code_0_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf10), .D(_22__1_), .Q(cond_code_1_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf9), .D(_22__2_), .Q(cond_code_2_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf10), .D(_30_), .Q(plp) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf10), .D(_29_), .Q(php) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf1), .D(_17_), .Q(clc) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf3), .D(_33_), .Q(sec) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf1), .D(_18_), .Q(cld) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf1), .D(_34_), .Q(sed) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf1), .D(_19_), .Q(cli) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf1), .D(_35_), .Q(sei) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf10), .D(_20_), .Q(clv) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf3), .D(_16_), .Q(bit_ins) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf3), .D(_28__0_), .Q(op_0_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf3), .D(_28__1_), .Q(op_1_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf3), .D(_28__2_), .Q(op_2_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf3), .D(_28__3_), .Q(op_3_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf1), .D(_32_), .Q(rotate) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf3), .D(_37_), .Q(shift_right) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf1), .D(_21_), .Q(compare) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf10), .D(_36_), .Q(shift) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf6), .D(_12_), .Q(adc_bcd) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf6), .D(_13_), .Q(adc_sbc) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf1), .D(_24_), .Q(inc) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf3), .D(_26_), .Q(load_only) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf10), .D(_40_), .Q(write_back) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf10), .D(_39_), .Q(store) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(new_wire_11), .D(_25_), .Q(index_y) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(new_wire_11), .D(_38__0_), .Q(src_reg_0_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(new_wire_20), .D(_38__1_), .Q(src_reg_1_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf9), .D(_23__0_), .Q(dst_reg_0_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(new_wire_11), .D(_23__1_), .Q(dst_reg_1_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(new_wire_11), .D(_27_), .Q(load_reg) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf4), .D(_31_), .Q(res) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf2), .D(DIMUX_0_), .Q(DIHOLD_0_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf4), .D(DIMUX_1_), .Q(DIHOLD_1_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf7), .D(DIMUX_2_), .Q(DIHOLD_2_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf2), .D(DIMUX_3_), .Q(DIHOLD_3_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf7), .D(DIMUX_4_), .Q(DIHOLD_4_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf2), .D(DIMUX_5_), .Q(DIHOLD_5_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf9), .D(DIMUX_6_), .Q(DIHOLD_6_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf9), .D(DIMUX_7_), .Q(DIHOLD_7_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf6), .D(_4__0_), .Q(IRHOLD_0_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf6), .D(_4__1_), .Q(IRHOLD_1_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf9), .D(_4__2_), .Q(IRHOLD_2_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf6), .D(_4__3_), .Q(IRHOLD_3_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf6), .D(_4__4_), .Q(IRHOLD_4_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf6), .D(_4__5_), .Q(IRHOLD_5_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf9), .D(_4__6_), .Q(IRHOLD_6_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(new_wire_20), .D(_4__7_), .Q(IRHOLD_7_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(new_wire_15), .D(_5_), .Q(IRHOLD_valid) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf9), .D(_10_), .Q(V) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf9), .D(_3_), .Q(D) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf7), .D(_6_), .Q(I) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(new_wire_12), .D(_8_), .Q(N) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(new_wire_12), .D(_11_), .Q(Z) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(new_wire_12), .D(_2_), .Q(C) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(new_wire_12), .D(_15_), .Q(backwards) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(new_wire_15), .D(_14_), .Q(adj_bcd) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf2), .D(_1__0_), .Q(ABL_0_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf0), .D(_1__1_), .Q(ABL_1_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf2), .D(_1__2_), .Q(ABL_2_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf2), .D(_1__3_), .Q(ABL_3_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf2), .D(_1__4_), .Q(ABL_4_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf2), .D(_1__5_), .Q(ABL_5_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(new_wire_10), .D(_1__6_), .Q(ABL_6_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(new_wire_19), .D(_1__7_), .Q(ABL_7_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf7), .D(_0__0_), .Q(ABH_0_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf0), .D(_0__1_), .Q(ABH_1_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(new_wire_19), .D(_0__2_), .Q(ABH_2_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf7), .D(_0__3_), .Q(ABH_3_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(new_wire_14), .D(_0__4_), .Q(ABH_4_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(new_wire_14), .D(_0__5_), .Q(ABH_5_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(new_wire_14), .D(_0__6_), .Q(ABH_6_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(new_wire_14), .D(_0__7_), .Q(ABH_7_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf4), .D(_9__0_), .Q(PC_0_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf0), .D(_9__1_), .Q(PC_1_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf0), .D(_9__2_), .Q(PC_2_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf0), .D(_9__3_), .Q(PC_3_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(new_wire_19), .D(_9__4_), .Q(PC_4_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf0), .D(_9__5_), .Q(PC_5_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf4), .D(_9__6_), .Q(PC_6_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf4), .D(_9__7_), .Q(PC_7_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf0), .D(_9__8_), .Q(PC_8_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf0), .D(_9__9_), .Q(PC_9_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(new_wire_21), .D(_9__10_), .Q(PC_10_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(new_wire_19), .D(_9__11_), .Q(PC_11_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(new_wire_21), .D(_9__12_), .Q(PC_12_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(new_wire_21), .D(_9__13_), .Q(PC_13_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf4), .D(_9__14_), .Q(PC_14_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(new_wire_21), .D(_9__15_), .Q(PC_15_) );
DFFSR DFFSR_1 ( .CLK(clk_bF_buf4), .D(_1438__0_), .Q(state_0_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_2 ( .CLK(clk_bF_buf4), .D(_1438__1_), .Q(state_1_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_3 ( .CLK(new_wire_17), .D(_1438__2_), .Q(state_2_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_4 ( .CLK(new_wire_17), .D(_1438__3_), .Q(state_3_), .R(vdd), .S(_1175_) );
DFFSR DFFSR_5 ( .CLK(new_wire_17), .D(_1438__4_), .Q(state_4_), .R(_1175_), .S(vdd) );
DFFSR DFFSR_6 ( .CLK(new_wire_17), .D(_1438__5_), .Q(state_5_), .R(_1175_), .S(vdd) );
OR2X2 OR2X2_38 ( .A(new_wire_50), .B(new_wire_49), .Y(_1626_) );
NOR2X1 NOR2X1_224 ( .A(new_wire_48), .B(new_wire_47), .Y(_1627_) );
NOR2X1 NOR2X1_225 ( .A(new_wire_45), .B(ADD_5_), .Y(_1628_) );
NOR2X1 NOR2X1_226 ( .A(new_wire_51), .B(ADD_1_), .Y(_1629_) );
NAND3X1 NAND3X1_164 ( .A(_1627_), .B(_1628_), .C(_1629_), .Y(_1630_) );
NOR2X1 NOR2X1_227 ( .A(_1626_), .B(_1630_), .Y(AZ) );
INVX8 INVX8_7 ( .A(new_wire_4), .Y(_1631_) );
NAND2X1 NAND2X1_212 ( .A(CO), .B(_1631__bF_buf3), .Y(_1632_) );
NOR2X1 NOR2X1_228 ( .A(alu_op_2_), .B(_1633_), .Y(_1634_) );
NOR2X1 NOR2X1_229 ( .A(alu_op_1_), .B(_1635_), .Y(_1636_) );
NOR2X1 NOR2X1_230 ( .A(alu_op_0_), .B(_1637_), .Y(_1638_) );
OAI21X1 OAI21X1_395 ( .A(_1639_), .B(_1640_), .C(BI_5_), .Y(_1641_) );
OAI21X1 OAI21X1_396 ( .A(_1636_), .B(_1638_), .C(_1641_), .Y(_1642_) );
AOI21X1 AOI21X1_121 ( .A(_1643_), .B(_1640_), .C(alu_shift_right), .Y(_1644_) );
AOI22X1 AOI22X1_51 ( .A(alu_shift_right), .B(AI_6_), .C(_1642_), .D(_1644_), .Y(_1645_) );
NOR2X1 NOR2X1_231 ( .A(alu_op_3_), .B(_1647_), .Y(_1648_) );
OAI21X1 OAI21X1_397 ( .A(alu_op_2_), .B(alu_op_3_), .C(BI_5_), .Y(_1649_) );
OAI21X1 OAI21X1_398 ( .A(BI_5_), .B(_1648_), .C(_1649_), .Y(_1650_) );
OAI21X1 OAI21X1_399 ( .A(_1634_), .B(_1651_), .C(_1646_), .Y(_1652_) );
NAND2X1 NAND2X1_213 ( .A(alu_op_0_), .B(_1639_), .Y(_1655_) );
AND2X2 AND2X2_48 ( .A(_1635_), .B(BI_4_), .Y(_1656_) );
NAND2X1 NAND2X1_214 ( .A(AI_4_), .B(_1656_), .Y(_1657_) );
AOI22X1 AOI22X1_52 ( .A(_1639_), .B(BI_4_), .C(_1655_), .D(_1657_), .Y(_1658_) );
OAI21X1 OAI21X1_400 ( .A(AI_4_), .B(_1656_), .C(_1654_), .Y(_1659_) );
OAI22X1 OAI22X1_55 ( .A(_1654_), .B(_1640_), .C(_1659_), .D(_1658_), .Y(_1660_) );
OAI21X1 OAI21X1_401 ( .A(alu_op_2_), .B(alu_op_3_), .C(BI_4_), .Y(_1661_) );
OAI21X1 OAI21X1_402 ( .A(BI_4_), .B(_1648_), .C(_1661_), .Y(_1662_) );
OAI21X1 OAI21X1_403 ( .A(_1634_), .B(_1663_), .C(_1660_), .Y(_1664_) );
NOR2X1 NOR2X1_232 ( .A(alu_op_0_), .B(_1666_), .Y(_1667_) );
OAI21X1 OAI21X1_404 ( .A(_1639_), .B(_1668_), .C(BI_2_), .Y(_1669_) );
OAI21X1 OAI21X1_405 ( .A(_1636_), .B(_1667_), .C(_1669_), .Y(_1670_) );
OAI21X1 OAI21X1_406 ( .A(alu_op_0_), .B(_1666_), .C(_1668_), .Y(_1671_) );
NAND3X1 NAND3X1_165 ( .A(_1654_), .B(_1671_), .C(_1670_), .Y(_1452_) );
OAI21X1 OAI21X1_407 ( .A(_1654_), .B(_1665_), .C(_1452_), .Y(_1453_) );
OAI21X1 OAI21X1_408 ( .A(alu_op_2_), .B(alu_op_3_), .C(BI_2_), .Y(_1454_) );
OAI21X1 OAI21X1_409 ( .A(BI_2_), .B(_1648_), .C(_1454_), .Y(_1455_) );
OAI21X1 OAI21X1_410 ( .A(alu_op_2_), .B(_1633_), .C(_1455_), .Y(_1456_) );
NAND3X1 NAND3X1_166 ( .A(AI_1_), .B(BI_1_), .C(_1635_), .Y(_1457_) );
AOI22X1 AOI22X1_53 ( .A(_1639_), .B(BI_1_), .C(_1655_), .D(_1457_), .Y(_1458_) );
OAI21X1 OAI21X1_411 ( .A(alu_op_0_), .B(_1460_), .C(_1459_), .Y(_1461_) );
NAND2X1 NAND2X1_215 ( .A(_1654_), .B(_1461_), .Y(_1462_) );
OAI22X1 OAI22X1_56 ( .A(_1654_), .B(_1668_), .C(_1462_), .D(_1458_), .Y(_1463_) );
OAI21X1 OAI21X1_412 ( .A(alu_op_2_), .B(alu_op_3_), .C(BI_1_), .Y(_1464_) );
OAI21X1 OAI21X1_413 ( .A(BI_1_), .B(_1648_), .C(_1464_), .Y(_1465_) );
OAI21X1 OAI21X1_414 ( .A(_1634_), .B(_1466_), .C(_1463_), .Y(_1467_) );
NAND2X1 NAND2X1_216 ( .A(alu_shift_right), .B(AI_1_), .Y(_1468_) );
NAND2X1 NAND2X1_217 ( .A(BI_0_), .B(_1635_), .Y(_1469_) );
NAND2X1 NAND2X1_218 ( .A(alu_op_1_), .B(AI_0_), .Y(_1470_) );
AOI22X1 AOI22X1_54 ( .A(BI_0_), .B(_1470_), .C(_1655_), .D(_1469_), .Y(_1471_) );
OAI21X1 OAI21X1_415 ( .A(alu_op_0_), .B(_1473_), .C(_1472_), .Y(_1474_) );
NAND2X1 NAND2X1_219 ( .A(_1654_), .B(_1474_), .Y(_1475_) );
OAI21X1 OAI21X1_416 ( .A(_1471_), .B(_1475_), .C(_1468_), .Y(_1476_) );
OAI21X1 OAI21X1_417 ( .A(alu_op_2_), .B(alu_op_3_), .C(BI_0_), .Y(_1477_) );
OAI21X1 OAI21X1_418 ( .A(BI_0_), .B(_1648_), .C(_1477_), .Y(_1478_) );
OAI21X1 OAI21X1_419 ( .A(new_wire_65), .B(_1633_), .C(_1478_), .Y(_1479_) );
OAI21X1 OAI21X1_420 ( .A(_1647_), .B(_1633_), .C(CI), .Y(_1480_) );
NOR2X1 NOR2X1_233 ( .A(alu_shift_right), .B(_1480_), .Y(_1481_) );
MUX2X1 MUX2X1_35 ( .A(alu_op_1_), .B(_1473_), .S(alu_op_0_), .Y(_1482_) );
NAND2X1 NAND2X1_220 ( .A(BI_0_), .B(_1470_), .Y(_1483_) );
NAND2X1 NAND2X1_221 ( .A(_1483_), .B(_1482_), .Y(_1484_) );
AOI21X1 AOI21X1_122 ( .A(_1469_), .B(_1472_), .C(alu_shift_right), .Y(_1485_) );
NAND2X1 NAND2X1_222 ( .A(_1485_), .B(_1484_), .Y(_1486_) );
NAND3X1 NAND3X1_167 ( .A(_1468_), .B(_1478_), .C(_1486_), .Y(_1487_) );
AOI22X1 AOI22X1_55 ( .A(_1476_), .B(_1479_), .C(_1481_), .D(_1487_), .Y(_1488_) );
NOR2X1 NOR2X1_234 ( .A(_1466_), .B(_1463_), .Y(_1489_) );
OAI21X1 OAI21X1_421 ( .A(_1489_), .B(_1488_), .C(_1467_), .Y(_1490_) );
MUX2X1 MUX2X1_36 ( .A(_1456_), .B(_1455_), .S(_1453_), .Y(_1491_) );
AOI22X1 AOI22X1_56 ( .A(_1453_), .B(_1456_), .C(_1491_), .D(_1490_), .Y(_1492_) );
NAND2X1 NAND2X1_223 ( .A(alu_shift_right), .B(AI_4_), .Y(_1493_) );
NOR2X1 NOR2X1_235 ( .A(new_wire_64), .B(_1494_), .Y(_1495_) );
NAND2X1 NAND2X1_224 ( .A(AI_3_), .B(_1495_), .Y(_1496_) );
AOI22X1 AOI22X1_57 ( .A(_1639_), .B(BI_3_), .C(_1655_), .D(_1496_), .Y(_1497_) );
OAI21X1 OAI21X1_422 ( .A(AI_3_), .B(_1495_), .C(_1654_), .Y(_1498_) );
OAI21X1 OAI21X1_423 ( .A(_1498_), .B(_1497_), .C(_1493_), .Y(_1499_) );
OAI21X1 OAI21X1_424 ( .A(alu_op_3_), .B(_1647_), .C(_1494_), .Y(_1500_) );
OAI21X1 OAI21X1_425 ( .A(new_wire_65), .B(new_wire_66), .C(BI_3_), .Y(_1501_) );
AND2X2 AND2X2_49 ( .A(_1500_), .B(_1501_), .Y(_1502_) );
OAI21X1 OAI21X1_426 ( .A(_1634_), .B(_1502_), .C(_1499_), .Y(_1503_) );
OAI21X1 OAI21X1_427 ( .A(_1499_), .B(_1502_), .C(_1503_), .Y(_1504_) );
XOR2X1 XOR2X1_2 ( .A(_1492_), .B(_1504_), .Y(_1505_) );
OAI21X1 OAI21X1_428 ( .A(_1634_), .B(_1507_), .C(_1476_), .Y(_1508_) );
NOR2X1 NOR2X1_236 ( .A(_1507_), .B(_1476_), .Y(_1510_) );
OAI21X1 OAI21X1_429 ( .A(_1509_), .B(_1510_), .C(_1508_), .Y(_1511_) );
OAI21X1 OAI21X1_430 ( .A(new_wire_65), .B(_1633_), .C(_1465_), .Y(_1512_) );
AOI21X1 AOI21X1_123 ( .A(_1463_), .B(_1512_), .C(_1489_), .Y(_1513_) );
NAND2X1 NAND2X1_225 ( .A(_1513_), .B(_1511_), .Y(_1514_) );
OAI21X1 OAI21X1_431 ( .A(_1463_), .B(_1466_), .C(_1467_), .Y(_1515_) );
NAND2X1 NAND2X1_226 ( .A(_1488_), .B(_1515_), .Y(_1516_) );
NAND2X1 NAND2X1_227 ( .A(_1516_), .B(_1514_), .Y(_1517_) );
NAND2X1 NAND2X1_228 ( .A(_1491_), .B(_1490_), .Y(_1518_) );
OAI21X1 OAI21X1_432 ( .A(_1634_), .B(_1519_), .C(_1453_), .Y(_1520_) );
OAI21X1 OAI21X1_433 ( .A(_1453_), .B(_1519_), .C(_1520_), .Y(_1521_) );
NAND3X1 NAND3X1_168 ( .A(_1467_), .B(_1521_), .C(_1514_), .Y(_1522_) );
NAND2X1 NAND2X1_229 ( .A(_1518_), .B(_1522_), .Y(_1523_) );
AOI21X1 AOI21X1_124 ( .A(_1523_), .B(_1517_), .C(_1506_), .Y(_1524_) );
OAI21X1 OAI21X1_434 ( .A(_1504_), .B(_1492_), .C(_1503_), .Y(_1525_) );
AOI21X1 AOI21X1_125 ( .A(_1524_), .B(_1505_), .C(_1525_), .Y(_1526_) );
OAI21X1 OAI21X1_435 ( .A(_1660_), .B(_1663_), .C(_1664_), .Y(_1527_) );
OAI21X1 OAI21X1_436 ( .A(_1527_), .B(_1526_), .C(_1664_), .Y(_1528_) );
OAI21X1 OAI21X1_437 ( .A(_1646_), .B(_1651_), .C(_1652_), .Y(_1529_) );
AOI21X1 AOI21X1_126 ( .A(_1528_), .B(_1530_), .C(_1653_), .Y(_1531_) );
NOR2X1 NOR2X1_237 ( .A(new_wire_64), .B(_1532_), .Y(_1533_) );
OAI21X1 OAI21X1_438 ( .A(_1639_), .B(_1534_), .C(BI_7_), .Y(_1535_) );
OAI21X1 OAI21X1_439 ( .A(_1636_), .B(_1533_), .C(_1535_), .Y(_1536_) );
AOI21X1 AOI21X1_127 ( .A(_1537_), .B(_1534_), .C(alu_shift_right), .Y(_1538_) );
AOI22X1 AOI22X1_58 ( .A(CI), .B(new_wire_70), .C(_1536_), .D(_1538_), .Y(_1539_) );
OAI21X1 OAI21X1_440 ( .A(new_wire_65), .B(new_wire_66), .C(BI_7_), .Y(_1541_) );
OAI21X1 OAI21X1_441 ( .A(BI_7_), .B(_1648_), .C(_1541_), .Y(_1542_) );
OAI21X1 OAI21X1_442 ( .A(_1543_), .B(_1634_), .C(_1540_), .Y(_1544_) );
NOR2X1 NOR2X1_238 ( .A(new_wire_64), .B(_1546_), .Y(_1547_) );
OAI21X1 OAI21X1_443 ( .A(_1639_), .B(_1548_), .C(BI_6_), .Y(_1549_) );
OAI21X1 OAI21X1_444 ( .A(_1636_), .B(_1547_), .C(_1549_), .Y(_1550_) );
AOI21X1 AOI21X1_128 ( .A(_1551_), .B(_1548_), .C(new_wire_70), .Y(_1552_) );
AOI22X1 AOI22X1_59 ( .A(AI_7_), .B(new_wire_70), .C(_1550_), .D(_1552_), .Y(_1553_) );
OAI21X1 OAI21X1_445 ( .A(new_wire_65), .B(new_wire_66), .C(BI_6_), .Y(_1555_) );
OAI21X1 OAI21X1_446 ( .A(BI_6_), .B(_1648_), .C(_1555_), .Y(_1556_) );
OAI21X1 OAI21X1_447 ( .A(_1634_), .B(_1557_), .C(_1554_), .Y(_1558_) );
OAI21X1 OAI21X1_448 ( .A(_1540_), .B(_1543_), .C(_1544_), .Y(_1560_) );
AOI21X1 AOI21X1_129 ( .A(_1561_), .B(_1559_), .C(_1545_), .Y(_1562_) );
OAI21X1 OAI21X1_449 ( .A(_1554_), .B(_1557_), .C(_1558_), .Y(_1563_) );
NAND2X1 NAND2X1_230 ( .A(_1564_), .B(_1561_), .Y(_1565_) );
OAI21X1 OAI21X1_450 ( .A(_1565_), .B(_1531_), .C(_1562_), .Y(_1566_) );
NAND3X1 NAND3X1_169 ( .A(new_wire_70), .B(AI_0_), .C(_1566_), .Y(_1567_) );
NAND2X1 NAND2X1_231 ( .A(new_wire_70), .B(AI_0_), .Y(_1568_) );
OR2X2 OR2X2_39 ( .A(_1531_), .B(_1565_), .Y(_1569_) );
NAND3X1 NAND3X1_170 ( .A(_1568_), .B(_1562_), .C(_1569_), .Y(_1570_) );
NAND2X1 NAND2X1_232 ( .A(_1505_), .B(_1524_), .Y(_1572_) );
OAI21X1 OAI21X1_451 ( .A(_1575_), .B(_1574_), .C(_1662_), .Y(_1576_) );
OR2X2 OR2X2_40 ( .A(_1576_), .B(_1574_), .Y(_1577_) );
NAND2X1 NAND2X1_233 ( .A(_1574_), .B(_1576_), .Y(_1578_) );
AOI22X1 AOI22X1_60 ( .A(_1577_), .B(_1578_), .C(_1573_), .D(_1572_), .Y(_1579_) );
OAI21X1 OAI21X1_452 ( .A(_1571_), .B(_1579_), .C(_1530_), .Y(_1580_) );
OAI21X1 OAI21X1_453 ( .A(_1575_), .B(_1553_), .C(_1556_), .Y(_1581_) );
OR2X2 OR2X2_41 ( .A(_1581_), .B(_1553_), .Y(_1582_) );
NAND2X1 NAND2X1_234 ( .A(_1553_), .B(_1581_), .Y(_1583_) );
AOI22X1 AOI22X1_61 ( .A(_1582_), .B(_1583_), .C(_1652_), .D(_1580_), .Y(_1584_) );
OAI21X1 OAI21X1_454 ( .A(_1559_), .B(_1584_), .C(_1560_), .Y(_1585_) );
OAI21X1 OAI21X1_455 ( .A(new_wire_65), .B(_1633_), .C(_1662_), .Y(_1586_) );
XNOR2X1 XNOR2X1_8 ( .A(_1492_), .B(_1504_), .Y(_1587_) );
NAND3X1 NAND3X1_171 ( .A(_1467_), .B(_1491_), .C(_1514_), .Y(_1588_) );
NAND2X1 NAND2X1_235 ( .A(_1521_), .B(_1490_), .Y(_1589_) );
NAND3X1 NAND3X1_172 ( .A(_1589_), .B(_1517_), .C(_1588_), .Y(_1590_) );
NAND2X1 NAND2X1_236 ( .A(ALU_BCD), .B(_1590_), .Y(_1591_) );
OAI21X1 OAI21X1_456 ( .A(_1591_), .B(_1587_), .C(_1573_), .Y(_1592_) );
AOI22X1 AOI22X1_62 ( .A(_1660_), .B(_1586_), .C(_1593_), .D(_1592_), .Y(_1594_) );
OAI21X1 OAI21X1_457 ( .A(_1529_), .B(_1594_), .C(_1652_), .Y(_1595_) );
NAND2X1 NAND2X1_237 ( .A(_1564_), .B(_1595_), .Y(_1596_) );
NAND3X1 NAND3X1_173 ( .A(_1558_), .B(_1561_), .C(_1596_), .Y(_1597_) );
NAND2X1 NAND2X1_238 ( .A(_1597_), .B(_1585_), .Y(_1598_) );
NAND2X1 NAND2X1_239 ( .A(_1529_), .B(_1594_), .Y(_1599_) );
NAND2X1 NAND2X1_240 ( .A(_1599_), .B(_1580_), .Y(_1600_) );
NAND3X1 NAND3X1_174 ( .A(_1652_), .B(_1563_), .C(_1580_), .Y(_1601_) );
NAND2X1 NAND2X1_241 ( .A(_1601_), .B(_1596_), .Y(_1602_) );
AOI21X1 AOI21X1_130 ( .A(_1602_), .B(_1600_), .C(_1506_), .Y(_1603_) );
AOI22X1 AOI22X1_63 ( .A(_1567_), .B(_1570_), .C(_1598_), .D(_1603_), .Y(_1604_) );
OAI21X1 OAI21X1_458 ( .A(_1631__bF_buf3), .B(_1604_), .C(_1632_), .Y(_1448_) );
NAND2X1 NAND2X1_242 ( .A(AN), .B(_1631__bF_buf2), .Y(_1606_) );
OAI21X1 OAI21X1_459 ( .A(_1631__bF_buf2), .B(_1605_), .C(_1606_), .Y(_1450_) );
NAND2X1 NAND2X1_243 ( .A(HC), .B(_1631__bF_buf0), .Y(_1607_) );
OAI21X1 OAI21X1_460 ( .A(_1631__bF_buf0), .B(_1526_), .C(_1607_), .Y(_1449_) );
NAND2X1 NAND2X1_244 ( .A(new_wire_49), .B(_1631__bF_buf1), .Y(_1608_) );
AOI21X1 AOI21X1_131 ( .A(_1508_), .B(_1487_), .C(_1481_), .Y(_1609_) );
OAI21X1 OAI21X1_461 ( .A(_1476_), .B(_1507_), .C(_1508_), .Y(_1610_) );
OAI21X1 OAI21X1_462 ( .A(_1509_), .B(_1610_), .C(new_wire_4), .Y(_1611_) );
OAI21X1 OAI21X1_463 ( .A(_1609_), .B(_1611_), .C(_1608_), .Y(_1451__0_) );
NAND2X1 NAND2X1_245 ( .A(ADD_1_), .B(_1631__bF_buf0), .Y(_1612_) );
OAI21X1 OAI21X1_464 ( .A(_1631__bF_buf0), .B(_1517_), .C(_1612_), .Y(_1451__1_) );
NAND2X1 NAND2X1_246 ( .A(new_wire_51), .B(_1631__bF_buf1), .Y(_1613_) );
OAI21X1 OAI21X1_465 ( .A(_1631__bF_buf1), .B(_1523_), .C(_1613_), .Y(_1451__2_) );
NAND2X1 NAND2X1_247 ( .A(new_wire_50), .B(_1631__bF_buf1), .Y(_1614_) );
OAI21X1 OAI21X1_466 ( .A(_1631__bF_buf1), .B(_1587_), .C(_1614_), .Y(_1451__3_) );
NAND2X1 NAND2X1_248 ( .A(new_wire_45), .B(_1631__bF_buf1), .Y(_1615_) );
NOR2X1 NOR2X1_239 ( .A(_1593_), .B(_1592_), .Y(_1616_) );
OAI21X1 OAI21X1_467 ( .A(_1527_), .B(_1526_), .C(new_wire_4), .Y(_1617_) );
OAI21X1 OAI21X1_468 ( .A(_1616_), .B(_1617_), .C(_1615_), .Y(_1451__4_) );
NAND2X1 NAND2X1_249 ( .A(new_wire_42), .B(_1631__bF_buf0), .Y(_1618_) );
OAI21X1 OAI21X1_469 ( .A(_1631__bF_buf0), .B(_1600_), .C(_1618_), .Y(_1451__5_) );
NAND2X1 NAND2X1_250 ( .A(new_wire_48), .B(_1631__bF_buf3), .Y(_1619_) );
OAI21X1 OAI21X1_470 ( .A(_1631__bF_buf3), .B(_1602_), .C(_1619_), .Y(_1451__6_) );
NAND2X1 NAND2X1_251 ( .A(new_wire_47), .B(_1631__bF_buf3), .Y(_1620_) );
OAI21X1 OAI21X1_471 ( .A(_1631__bF_buf3), .B(_1605_), .C(_1620_), .Y(_1451__7_) );
AOI21X1 AOI21X1_132 ( .A(_1540_), .B(new_wire_79), .C(_1543_), .Y(_1621_) );
NAND2X1 NAND2X1_252 ( .A(ALU_BI7), .B(_1631__bF_buf2), .Y(_1622_) );
OAI21X1 OAI21X1_472 ( .A(_1631__bF_buf2), .B(_1621_), .C(_1622_), .Y(_1447_) );
NAND2X1 NAND2X1_253 ( .A(ALU_AI7), .B(_1631__bF_buf2), .Y(_1623_) );
OAI21X1 OAI21X1_473 ( .A(_1534_), .B(_1631__bF_buf2), .C(_1623_), .Y(_1446_) );
XOR2X1 XOR2X1_3 ( .A(ALU_BI7), .B(ALU_AI7), .Y(_1624_) );
XNOR2X1 XNOR2X1_9 ( .A(CO), .B(AN), .Y(_1625_) );
XNOR2X1 XNOR2X1_10 ( .A(_1624_), .B(_1625_), .Y(AV) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(new_wire_20), .D(_1448_), .Q(CO) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(new_wire_18), .D(_1450_), .Q(AN) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(new_wire_15), .D(_1449_), .Q(HC) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(new_wire_13), .D(_1451__0_), .Q(ADD_0_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(new_wire_16), .D(_1451__1_), .Q(ADD_1_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(new_wire_13), .D(_1451__2_), .Q(ADD_2_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(new_wire_16), .D(_1451__3_), .Q(ADD_3_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(new_wire_16), .D(_1451__4_), .Q(ADD_4_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(new_wire_15), .D(_1451__5_), .Q(ADD_5_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(new_wire_18), .D(_1451__6_), .Q(ADD_6_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(new_wire_20), .D(_1451__7_), .Q(ADD_7_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(new_wire_18), .D(_1447_), .Q(ALU_BI7) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(new_wire_18), .D(_1446_), .Q(ALU_AI7) );
BUFX4 BUFX4_1_clone_[1] ( .A(RDY), .Y(new_wire_1) );
BUFX4 BUFX4_2_clone_[2] ( .A(RDY), .Y(new_wire_2) );
BUFX4 BUFX4_3_clone_[3] ( .A(RDY), .Y(new_wire_3) );
BUFX4 BUFX4_4_clone_[4] ( .A(RDY), .Y(new_wire_4) );
BUFX4 BUFX4_5_clone_[5] ( .A(RDY), .Y(new_wire_5) );
BUFX4 BUFX4_6_clone_[6] ( .A(RDY), .Y(new_wire_6) );
BUFX4 BUFX4_7_clone_[7] ( .A(RDY), .Y(new_wire_7) );
BUFX4 BUFX4_8_clone_[8] ( .A(RDY), .Y(new_wire_8) );
BUFX4 BUFX4_9_clone_[9] ( .A(RDY), .Y(new_wire_9) );
BUFX4 BUFX4_15_clone_[10] ( .A(clk), .Y(new_wire_10) );
BUFX4 BUFX4_16_clone_[11] ( .A(clk), .Y(new_wire_11) );
BUFX4 BUFX4_17_clone_[12] ( .A(clk), .Y(new_wire_12) );
BUFX4 BUFX4_18_clone_[13] ( .A(clk), .Y(new_wire_13) );
BUFX4 BUFX4_19_clone_[14] ( .A(clk), .Y(new_wire_14) );
BUFX4 BUFX4_20_clone_[15] ( .A(clk), .Y(new_wire_15) );
BUFX4 BUFX4_21_clone_[16] ( .A(clk), .Y(new_wire_16) );
BUFX4 BUFX4_22_clone_[17] ( .A(clk), .Y(new_wire_17) );
BUFX4 BUFX4_23_clone_[18] ( .A(clk), .Y(new_wire_18) );
BUFX4 BUFX4_24_clone_[19] ( .A(clk), .Y(new_wire_19) );
BUFX4 BUFX4_25_clone_[20] ( .A(clk), .Y(new_wire_20) );
BUFX4 BUFX4_26_clone_[21] ( .A(clk), .Y(new_wire_21) );
BUFX4 BUFX4_67_clone_[22] ( .A(new_wire_23), .Y(new_wire_22) );
INVX8 INVX8_5_clone_[23] ( .A(new_wire_24), .Y(new_wire_23) );
BUFX4 BUFX4_7_clone_[24] ( .A(RDY), .Y(new_wire_24) );
BUFX4 BUFX4_68_clone_[25] ( .A(new_wire_26), .Y(new_wire_25) );
INVX8 INVX8_5_clone_[26] ( .A(new_wire_27), .Y(new_wire_26) );
BUFX4 BUFX4_7_clone_[27] ( .A(RDY), .Y(new_wire_27) );
BUFX4 BUFX4_69_clone_[28] ( .A(new_wire_29), .Y(new_wire_28) );
INVX8 INVX8_5_clone_[29] ( .A(new_wire_30), .Y(new_wire_29) );
BUFX4 BUFX4_7_clone_[30] ( .A(RDY), .Y(new_wire_30) );
NOR2X1 NOR2X1_2_clone_[31] ( .A(state_5_), .B(_793_), .Y(new_wire_31) );
NOR2X1 NOR2X1_4_clone_[32] ( .A(state_4_), .B(_797_), .Y(new_wire_32) );
NOR2X1 NOR2X1_7_clone_[33] ( .A(_796_), .B(_807_), .Y(new_wire_33) );
NAND3X1 NAND3X1_2_clone_[34] ( .A(_812__bF_buf1), .B(_805_), .C(_814_), .Y(new_wire_34) );
NOR2X1 NOR2X1_11_clone_[35] ( .A(_816_), .B(_818_), .Y(new_wire_35) );
NAND2X1 NAND2X1_6_clone_[36] ( .A(new_wire_37), .B(new_wire_39), .Y(new_wire_36) );
NOR2X1 NOR2X1_7_clone_[37] ( .A(new_wire_38), .B(_807_), .Y(new_wire_37) );
NOR2X1 NOR2X1_3_clone_[38] ( .A(_795__bF_buf2), .B(_792_), .Y(new_wire_38) );
NOR2X1 NOR2X1_11_clone_[39] ( .A(_816_), .B(_818_), .Y(new_wire_39) );
INVX8 INVX8_3_clone_[40] ( .A(NMI_edge), .Y(new_wire_40) );
NAND3X1 NAND3X1_4_clone_[41] ( .A(_835_), .B(_839_), .C(_842_), .Y(new_wire_41) );
DFFPOSX1 DFFPOSX1_134_clone_[42] ( .CLK(new_wire_15), .D(_1451__5_), .Q(new_wire_42) );
NOR3X1 NOR3X1_2_clone_[43] ( .A(_809__bF_buf4), .B(_840_), .C(_848_), .Y(new_wire_43) );
NAND2X1 NAND2X1_16_clone_[44] ( .A(IRQ), .B(_828_), .Y(new_wire_44) );
DFFPOSX1 DFFPOSX1_133_clone_[45] ( .CLK(new_wire_16), .D(_1451__4_), .Q(new_wire_45) );
DFFPOSX1 DFFPOSX1_136_clone_[47] ( .CLK(new_wire_20), .D(_1451__7_), .Q(new_wire_47) );
DFFPOSX1 DFFPOSX1_135_clone_[48] ( .CLK(new_wire_18), .D(_1451__6_), .Q(new_wire_48) );
DFFPOSX1 DFFPOSX1_129_clone_[49] ( .CLK(new_wire_13), .D(_1451__0_), .Q(new_wire_49) );
DFFPOSX1 DFFPOSX1_132_clone_[50] ( .CLK(new_wire_16), .D(_1451__3_), .Q(new_wire_50) );
DFFPOSX1 DFFPOSX1_131_clone_[51] ( .CLK(new_wire_13), .D(_1451__2_), .Q(new_wire_51) );
DFFPOSX1 DFFPOSX1_85_clone_[52] ( .CLK(new_wire_15), .D(_5_), .Q(new_wire_52) );
NAND2X1 NAND2X1_45_clone_[53] ( .A(_830__bF_buf0), .B(_1089_), .Y(new_wire_53) );
NOR2X1 NOR2X1_45_clone_[54] ( .A(_825__bF_buf0), .B(_1093_), .Y(new_wire_54) );
AND2X2 AND2X2_10_clone_[56] ( .A(_1092_), .B(_830__bF_buf2), .Y(new_wire_56) );
NAND2X1 NAND2X1_57_clone_[57] ( .A(_802_), .B(_814_), .Y(new_wire_57) );
NAND2X1 NAND2X1_70_clone_[58] ( .A(_830__bF_buf1), .B(_1092_), .Y(new_wire_58) );
NOR2X1 NOR2X1_88_clone_[59] ( .A(_795__bF_buf4), .B(new_wire_60), .Y(new_wire_59) );
NAND2X1 NAND2X1_67_clone_[60] ( .A(_805_), .B(_814_), .Y(new_wire_60) );
OAI21X1 OAI21X1_147_clone_[61] ( .A(_128_), .B(_140_), .C(_144_), .Y(new_wire_61) );
OAI21X1 OAI21X1_147_clone_[63] ( .A(_128_), .B(_140_), .C(_144_), .Y(new_wire_63) );
OAI21X1 OAI21X1_162_clone_[64] ( .A(_266_), .B(_267_), .C(_273_), .Y(new_wire_64) );
OAI21X1 OAI21X1_164_clone_[65] ( .A(_275_), .B(_815__bF_buf1), .C(_277_), .Y(new_wire_65) );
NOR2X1 NOR2X1_146_clone_[66] ( .A(_278_), .B(_267_), .Y(new_wire_66) );
OAI21X1 OAI21X1_165_clone_[67] ( .A(_799__bF_buf3), .B(new_wire_68), .C(_271_), .Y(new_wire_67) );
NAND2X1 NAND2X1_57_clone_[68] ( .A(_802_), .B(new_wire_69), .Y(new_wire_68) );
NOR2X1 NOR2X1_10_clone_[69] ( .A(state_0_), .B(_813_), .Y(new_wire_69) );
AND2X2 AND2X2_41_clone_[70] ( .A(_81_), .B(shift_right), .Y(new_wire_70) );
NAND2X1 NAND2X1_166_clone_[71] ( .A(new_wire_62), .B(_470_), .Y(new_wire_71) );
OR2X2 OR2X2_21_clone_[72] ( .A(_524_), .B(reset), .Y(new_wire_72) );
NAND2X1 NAND2X1_180_clone_[73] ( .A(new_wire_61), .B(_470_), .Y(new_wire_73) );
NOR2X1 NOR2X1_193_clone_[74] ( .A(_95_), .B(_270_), .Y(new_wire_74) );
NAND3X1 NAND3X1_149_clone_[75] ( .A(_603_), .B(_600_), .C(_595_), .Y(new_wire_75) );
OAI21X1 OAI21X1_310_clone_[76] ( .A(_799__bF_buf4), .B(_1138_), .C(_1320_), .Y(new_wire_76) );
OR2X2 OR2X2_25_clone_[77] ( .A(_612_), .B(new_wire_78), .Y(new_wire_77) );
NAND3X1 NAND3X1_149_clone_[78] ( .A(_603_), .B(_600_), .C(_595_), .Y(new_wire_78) );
NOR2X1 NOR2X1_228_clone_[79] ( .A(new_wire_80), .B(_1633_), .Y(new_wire_79) );
OAI21X1 OAI21X1_164_clone_[80] ( .A(_275_), .B(_815__bF_buf1), .C(_277_), .Y(new_wire_80) );
BUFX4 BUFX2_1_s ( .A(_155_), .Y(_155__bF_buf3) );
BUFX4 BUFX2_2_s ( .A(_155_), .Y(_155__bF_buf2) );
BUFX4 BUFX2_3_s ( .A(_155_), .Y(_155__bF_buf1) );
BUFX4 BUFX2_4_s ( .A(_155_), .Y(_155__bF_buf0) );
BUFX4 BUFX2_5_s ( .A(_152_), .Y(_152__bF_buf1) );
BUFX4 BUFX2_6_s ( .A(_152_), .Y(_152__bF_buf0) );
BUFX4 BUFX2_7_s ( .A(_830_), .Y(_830__bF_buf3) );
BUFX4 BUFX2_8_s ( .A(_830_), .Y(_830__bF_buf2) );
BUFX4 BUFX2_9_s ( .A(_830_), .Y(_830__bF_buf1) );
BUFX4 BUFX2_10_s ( .A(_830_), .Y(_830__bF_buf0) );
BUFX4 BUFX2_11_s ( .A(_859_), .Y(_859__bF_buf1) );
BUFX4 BUFX2_12_s ( .A(_859_), .Y(_859__bF_buf0) );
BUFX4 BUFX2_13_s ( .A(_148_), .Y(_148__bF_buf2) );
BUFX4 BUFX2_14_s ( .A(_148_), .Y(_148__bF_buf1) );
BUFX4 BUFX2_15_s ( .A(_148_), .Y(_148__bF_buf0) );
BUFX4 BUFX2_16_s ( .A(_812_), .Y(_812__bF_buf2) );
INVX4 INVX1_1_s_s_s_s ( .A(PC_13_), .Y(_787_) );
INVX2 INVX2_1_s_s ( .A(_788_), .Y(_789_) );
INVX2 INVX1_2_s_s_s ( .A(state_2_), .Y(_790_) );
INVX2 INVX1_3_s_s_s ( .A(state_4_), .Y(_793_) );
INVX2 INVX1_4_s_s_s ( .A(state_5_), .Y(_797_) );
INVX2 INVX1_5_s_s_s ( .A(state_0_), .Y(_800_) );
INVX2 INVX1_6_s_s_s ( .A(state_3_), .Y(_804_) );
INVX2 INVX1_7_s_s_s ( .A(state_1_), .Y(_813_) );
INVX2 INVX1_8_s_s_s ( .A(_820_), .Y(_821_) );
INVX8 INVX1_9_s_s_s ( .A(IRQ), .Y(_823_) );
INVX4 INVX2_2_s_s_s ( .A(I), .Y(_828_) );
INVX2 INVX1_10_s_s_s ( .A(DIHOLD_5_), .Y(_844_) );
INVX4 INVX2_3_s_s_s ( .A(ADD_5_), .Y(_846_) );
INVX4 INVX2_4_s_s_s ( .A(PC_5_), .Y(_860_) );
INVX4 INVX1_11_s_s_s_s ( .A(ABL_5_), .Y(_862_) );
INVX4 INVX4_1_s_s ( .A(_847_), .Y(_870_) );
INVX4 INVX2_5_s_s_s ( .A(PC_4_), .Y(_872_) );
INVX4 INVX1_12_s_s_s_s ( .A(ABL_4_), .Y(_874_) );
INVX4 INVX2_6_s_s_s ( .A(PC_7_), .Y(_883_) );
INVX4 INVX1_13_s_s_s_s ( .A(ABL_7_), .Y(_885_) );
INVX4 INVX2_7_s_s_s ( .A(PC_6_), .Y(_893_) );
INVX4 INVX1_14_s_s_s_s ( .A(ABL_6_), .Y(_895_) );
INVX4 INVX2_8_s_s_s ( .A(ADD_0_), .Y(_904_) );
INVX4 INVX2_9_s_s_s ( .A(PC_0_), .Y(_905_) );
INVX2 INVX1_15_s_s_s ( .A(_842_), .Y(_911_) );
INVX2 INVX1_16_s_s_s ( .A(_920_), .Y(_921_) );
INVX2 INVX2_10_s_s ( .A(_923_), .Y(_924_) );
INVX4 INVX2_11_s_s_s ( .A(ADD_1_), .Y(_931_) );
INVX4 INVX2_12_s_s_s ( .A(PC_1_), .Y(_933_) );
INVX4 INVX2_13_s_s_s ( .A(PC_3_), .Y(_944_) );
INVX4 INVX1_17_s_s_s_s ( .A(ABL_3_), .Y(_946_) );
INVX2 INVX1_18_s_s_s ( .A(_952_), .Y(_953_) );
INVX4 INVX2_14_s_s_s ( .A(PC_2_), .Y(_956_) );
INVX4 INVX1_19_s_s_s_s ( .A(ABL_2_), .Y(_958_) );
INVX2 INVX1_20_s_s_s ( .A(DIHOLD_3_), .Y(_966_) );
INVX4 INVX1_21_s_s_s_s ( .A(ABH_3_), .Y(_970_) );
INVX4 INVX2_15_s_s_s ( .A(PC_11_), .Y(_972_) );
INVX4 INVX2_16_s_s_s ( .A(_978_), .Y(DIMUX_2_) );
INVX4 INVX1_22_s_s_s_s ( .A(ABH_2_), .Y(_981_) );
INVX4 INVX2_17_s_s_s ( .A(PC_10_), .Y(_983_) );
INVX2 INVX1_23_s_s_s ( .A(DIHOLD_1_), .Y(_990_) );
INVX4 INVX1_24_s_s_s_s ( .A(ABH_1_), .Y(_994_) );
INVX4 INVX2_18_s_s_s ( .A(PC_9_), .Y(_996_) );
INVX2 INVX1_25_s_s_s ( .A(DIHOLD_0_), .Y(_1002_) );
INVX4 INVX1_26_s_s_s_s ( .A(ABH_0_), .Y(_1006_) );
INVX4 INVX2_19_s_s_s ( .A(PC_8_), .Y(_1008_) );
INVX4 INVX2_20_s_s_s ( .A(PC_12_), .Y(_1016_) );
INVX2 INVX2_21_s_s ( .A(_1019_), .Y(DIMUX_4_) );
INVX4 INVX2_22_s_s_s ( .A(ABH_4_), .Y(_1020_) );
INVX2 INVX1_27_s_s_s ( .A(_941_), .Y(_1032_) );
INVX2 INVX1_28_s_s_s ( .A(_951_), .Y(_1036_) );
INVX4 INVX1_29_s_s_s_s ( .A(ABH_6_), .Y(_1049_) );
INVX4 INVX2_23_s_s_s ( .A(_1052_), .Y(DIMUX_6_) );
INVX4 INVX1_30_s_s_s_s ( .A(PC_15_), .Y(_1059_) );
INVX4 INVX1_31_s_s_s_s ( .A(ABH_7_), .Y(_1061_) );
INVX4 INVX2_24_s_s_s ( .A(_1064_), .Y(DIMUX_7_) );
INVX1 INVX1_32_s_s ( .A(_1066_), .Y(_1067_) );
INVX8 INVX4_2_s ( .A(IRHOLD_valid), .Y(_1073_) );
INVX2 INVX1_33_s_s_s ( .A(IRHOLD_3_), .Y(_1074_) );
INVX4 INVX4_3_s_s ( .A(_1099_), .Y(_1100_) );
INVX2 INVX1_34_s_s_s ( .A(_914_), .Y(_1106_) );
INVX2 INVX1_35_s_s_s ( .A(_1110_), .Y(_1111_) );
INVX4 INVX2_25_s_s_s ( .A(_1137_), .Y(_1138_) );
INVX2 INVX1_36_s_s_s ( .A(_1143_), .Y(_1144_) );
INVX2 INVX1_37_s_s_s ( .A(_1152_), .Y(_1153_) );
INVX2 INVX1_38_s_s_s ( .A(_1168_), .Y(_1169_) );
INVX4 INVX2_26_s_s_s ( .A(DIMUX_3_), .Y(_1179_) );
INVX1 INVX1_39_s_s ( .A(_1145_), .Y(_1191_) );
INVX2 INVX1_40_s_s_s ( .A(_1201_), .Y(_1202_) );
INVX4 INVX1_41_s_s_s_s ( .A(write_back), .Y(_1212_) );
INVX2 INVX2_27_s_s ( .A(_1244_), .Y(_1245_) );
INVX1 INVX1_42_s_s ( .A(_1243_), .Y(_1258_) );
INVX2 INVX1_43_s_s_s ( .A(IRHOLD_0_), .Y(_1262_) );
INVX1 INVX1_44_s_s ( .A(_1292_), .Y(_1293_) );
INVX2 INVX1_45_s_s_s ( .A(_1160_), .Y(_1297_) );
INVX2 INVX1_46_s_s_s ( .A(Z), .Y(_1303_) );
INVX4 INVX2_28_s_s_s ( .A(V), .Y(_1306_) );
INVX2 INVX1_47_s_s_s ( .A(_1230_), .Y(_1312_) );
INVX2 INVX1_48_s_s_s ( .A(_915_), .Y(_1319_) );
INVX1 INVX1_49_s_s ( .A(_1333_), .Y(_1334_) );
INVX1 INVX1_50_s_s ( .A(_1205_), .Y(_1338_) );
INVX2 INVX1_51_s_s_s ( .A(_1196_), .Y(_1376_) );
INVX2 INVX1_52_s_s_s ( .A(_1378_), .Y(_1379_) );
INVX4 INVX2_29_s_s_s ( .A(_1358_), .Y(_1388_) );
INVX2 INVX1_53_s_s_s ( .A(_1197_), .Y(_1394_) );
INVX2 INVX1_54_s_s_s ( .A(_1127_), .Y(_1404_) );
INVX2 INVX1_55_s_s_s ( .A(_1409_), .Y(_1410_) );
INVX4 INVX2_30_s_s_s ( .A(_1291_), .Y(_43_) );
INVX2 INVX1_56_s_s_s ( .A(_1234_), .Y(_52_) );
INVX2 INVX1_57_s_s_s ( .A(_1325_), .Y(_63_) );
INVX2 INVX1_58_s_s_s ( .A(_1272_), .Y(_65_) );
INVX2 INVX1_59_s_s_s ( .A(_1418_), .Y(_71_) );
INVX4 INVX1_60_s_s_s_s ( .A(C), .Y(_79_) );
INVX2 INVX1_61_s_s_s ( .A(rotate), .Y(_85_) );
INVX4 INVX2_31_s_s_s ( .A(compare), .Y(_86_) );
INVX4 INVX2_32_s_s_s ( .A(shift), .Y(_87_) );
INVX2 INVX1_62_s_s_s ( .A(_80_), .Y(_88_) );
INVX2 INVX1_63_s_s_s ( .A(_1206_), .Y(_91_) );
INVX2 INVX1_64_s_s_s ( .A(_1251_), .Y(_97_) );
INVX2 INVX1_65_s_s_s ( .A(_98_), .Y(_99_) );
INVX4 INVX2_33_s_s_s ( .A(DIMUX_0_), .Y(_104_) );
INVX4 INVX2_34_s_s_s ( .A(_1323_), .Y(_114_) );
INVX4 INVX2_35_s_s_s ( .A(DIMUX_1_), .Y(_118_) );
INVX2 INVX1_66_s_s_s ( .A(DIMUX_5_), .Y(_119_) );
INVX4 INVX4_4_s_s ( .A(_124_), .Y(_125_) );
INVX4 INVX1_67_s_s_s_s ( .A(src_reg_1_), .Y(_128_) );
INVX2 INVX1_68_s_s_s ( .A(dst_reg_1_), .Y(_141_) );
INVX2 INVX1_69_s_s_s ( .A(_143_), .Y(_144_) );
INVX4 INVX4_5_s_s ( .A(_145_), .Y(_146_) );
INVX2 INVX1_70_s_s_s ( .A(AXYS_1__0_), .Y(_147_) );
INVX2 INVX1_71_s_s_s ( .A(AXYS_0__0_), .Y(_154_) );
INVX2 INVX1_72_s_s_s ( .A(AXYS_3__0_), .Y(_158_) );
INVX2 INVX1_73_s_s_s ( .A(AXYS_2__0_), .Y(_160_) );
INVX2 INVX1_74_s_s_s ( .A(_1392_), .Y(_169_) );
INVX2 INVX1_75_s_s_s ( .A(AXYS_1__1_), .Y(_176_) );
INVX2 INVX1_76_s_s_s ( .A(AXYS_0__1_), .Y(_178_) );
INVX2 INVX1_77_s_s_s ( .A(AXYS_3__1_), .Y(_181_) );
INVX2 INVX1_78_s_s_s ( .A(AXYS_2__1_), .Y(_183_) );
INVX2 INVX1_79_s_s_s ( .A(AXYS_1__2_), .Y(_189_) );
INVX2 INVX1_80_s_s_s ( .A(AXYS_0__2_), .Y(_191_) );
INVX2 INVX1_81_s_s_s ( .A(AXYS_3__2_), .Y(_194_) );
INVX2 INVX1_82_s_s_s ( .A(AXYS_2__2_), .Y(_196_) );
INVX2 INVX1_83_s_s_s ( .A(AXYS_1__3_), .Y(_202_) );
INVX2 INVX1_84_s_s_s ( .A(AXYS_0__3_), .Y(_204_) );
INVX2 INVX1_85_s_s_s ( .A(AXYS_3__3_), .Y(_207_) );
INVX2 INVX1_86_s_s_s ( .A(AXYS_2__3_), .Y(_209_) );
INVX2 INVX1_87_s_s_s ( .A(AXYS_1__4_), .Y(_215_) );
INVX2 INVX1_88_s_s_s ( .A(AXYS_0__4_), .Y(_217_) );
INVX2 INVX1_89_s_s_s ( .A(AXYS_3__4_), .Y(_220_) );
INVX2 INVX1_90_s_s_s ( .A(AXYS_2__4_), .Y(_222_) );
INVX4 INVX1_91_s_s_s_s ( .A(ABH_5_), .Y(_226_) );
INVX2 INVX1_92_s_s_s ( .A(AXYS_1__5_), .Y(_229_) );
INVX2 INVX1_93_s_s_s ( .A(AXYS_0__5_), .Y(_231_) );
INVX2 INVX1_94_s_s_s ( .A(AXYS_3__5_), .Y(_234_) );
INVX2 INVX1_95_s_s_s ( .A(AXYS_2__5_), .Y(_236_) );
INVX2 INVX1_96_s_s_s ( .A(AXYS_1__6_), .Y(_242_) );
INVX2 INVX1_97_s_s_s ( .A(AXYS_0__6_), .Y(_244_) );
INVX2 INVX1_98_s_s_s ( .A(AXYS_3__6_), .Y(_247_) );
INVX2 INVX1_99_s_s_s ( .A(AXYS_2__6_), .Y(_249_) );
INVX2 INVX1_100_s_s_s ( .A(AXYS_1__7_), .Y(_255_) );
INVX2 INVX1_101_s_s_s ( .A(AXYS_0__7_), .Y(_257_) );
INVX2 INVX1_102_s_s_s ( .A(AXYS_3__7_), .Y(_260_) );
INVX2 INVX1_103_s_s_s ( .A(AXYS_2__7_), .Y(_262_) );
INVX4 INVX1_104_s_s_s_s ( .A(op_0_), .Y(_266_) );
INVX4 INVX1_105_s_s_s_s ( .A(_81_), .Y(_267_) );
INVX4 INVX2_36_s_s_s ( .A(_132_), .Y(_269_) );
INVX2 INVX1_106_s_s_s ( .A(op_1_), .Y(_274_) );
INVX4 INVX1_107_s_s_s_s ( .A(backwards), .Y(_275_) );
INVX2 INVX1_108_s_s_s ( .A(_271_), .Y(_276_) );
INVX4 INVX1_109_s_s_s_s ( .A(op_3_), .Y(_278_) );
INVX2 INVX1_110_s_s_s ( .A(store), .Y(_279_) );
INVX1 INVX1_111_s_s ( .A(_280_), .Y(_281_) );
INVX4 INVX2_37_s_s_s ( .A(_1192_), .Y(_283_) );
INVX4 INVX2_38_s_s_s ( .A(_106_), .Y(_287_) );
INVX4 INVX1_112_s_s_s_s ( .A(php), .Y(_290_) );
INVX2 INVX1_113_s_s_s ( .A(_293_), .Y(_294_) );
INVX2 INVX1_114_s_s_s ( .A(_291_), .Y(_314_) );
INVX4 INVX1_115_s_s_s_s ( .A(N), .Y(_318_) );
INVX4 INVX1_116_s_s_s_s ( .A(adc_bcd), .Y(_322_) );
INVX8 INVX4_6_s ( .A(reset), .Y(_1175_) );
INVX2 INVX1_117_s_s_s ( .A(res), .Y(_323_) );
INVX4 INVX2_39_s_s_s ( .A(plp), .Y(_324_) );
INVX2 INVX1_118_s_s_s ( .A(_916_), .Y(_328_) );
INVX4 INVX2_40_s_s_s ( .A(_1155_), .Y(_330_) );
INVX2 INVX1_119_s_s_s ( .A(sei), .Y(_331_) );
INVX2 INVX1_120_s_s_s ( .A(load_reg), .Y(_338_) );
INVX2 INVX1_121_s_s_s ( .A(_349_), .Y(_350_) );
INVX1 INVX1_122_s_s ( .A(_355_), .Y(_356_) );
INVX4 INVX1_123_s_s_s_s ( .A(new_wire_51), .Y(_360_) );
INVX4 INVX2_41_s_s_s ( .A(ADD_3_), .Y(_363_) );
INVX4 INVX1_124_s_s_s_s ( .A(ADD_4_), .Y(_367_) );
INVX4 INVX1_125_s_s_s_s ( .A(CO), .Y(_370_) );
INVX2 INVX1_126_s_s_s ( .A(_373_), .Y(_374_) );
INVX1 INVX1_127_s_s ( .A(_379_), .Y(_380_) );
INVX4 INVX1_128_s_s_s_s ( .A(ADD_6_), .Y(_384_) );
INVX4 INVX2_42_s_s_s ( .A(ADD_7_), .Y(_387_) );
INVX2 INVX1_129_s_s_s ( .A(NMI_1), .Y(_391_) );
INVX2 INVX1_130_s_s_s ( .A(_1097_), .Y(_397_) );
INVX2 INVX1_131_s_s_s ( .A(_398_), .Y(_399_) );
INVX2 INVX1_132_s_s_s ( .A(_404_), .Y(_405_) );
INVX2 INVX1_133_s_s_s ( .A(_418_), .Y(_419_) );
INVX2 INVX1_134_s_s_s ( .A(_408_), .Y(_424_) );
INVX2 INVX1_135_s_s_s ( .A(_1183_), .Y(_425_) );
INVX1 INVX1_136_s_s ( .A(_436_), .Y(_437_) );
INVX2 INVX1_137_s_s_s ( .A(_441_), .Y(_442_) );
INVX2 INVX1_138_s_s_s ( .A(_435_), .Y(_444_) );
INVX2 INVX1_139_s_s_s ( .A(_461_), .Y(_462_) );
INVX4 INVX2_43_s_s_s ( .A(adc_sbc), .Y(_466_) );
INVX2 INVX1_140_s_s_s ( .A(_415_), .Y(_482_) );
INVX2 INVX1_141_s_s_s ( .A(src_reg_0_), .Y(_489_) );
INVX2 INVX1_142_s_s_s ( .A(_491_), .Y(_492_) );
INVX2 INVX1_143_s_s_s ( .A(_430_), .Y(_495_) );
INVX2 INVX1_144_s_s_s ( .A(dst_reg_0_), .Y(_506_) );
INVX2 INVX1_145_s_s_s ( .A(IRHOLD_4_), .Y(_530_) );
INVX2 INVX1_146_s_s_s ( .A(IRHOLD_5_), .Y(_531_) );
INVX2 INVX1_147_s_s_s ( .A(IRHOLD_6_), .Y(_532_) );
INVX2 INVX1_148_s_s_s ( .A(IRHOLD_7_), .Y(_533_) );
INVX4 INVX1_149_s_s_s_s ( .A(bit_ins), .Y(_539_) );
INVX4 INVX1_150_s_s_s_s ( .A(AN), .Y(_559_) );
INVX2 INVX1_151_s_s_s ( .A(AZ), .Y(_570_) );
INVX2 INVX1_152_s_s_s ( .A(ABL_0_), .Y(_614_) );
INVX2 INVX1_153_s_s_s ( .A(_135_), .Y(_621_) );
INVX2 INVX1_154_s_s_s ( .A(_142_), .Y(_647_) );
INVX2 INVX1_155_s_s_s ( .A(ABL_1_), .Y(_654_) );
INVX4 INVX2_44_s_s_s ( .A(_600_), .Y(_702_) );
INVX4 INVX4_7_s_s ( .A(_608_), .Y(_703_) );
INVX2 INVX1_156_s_s_s ( .A(PC_14_), .Y(_723_) );
INVX2 INVX1_157_s_s_s ( .A(_902_), .Y(_734_) );
INVX2 INVX1_158_s_s_s ( .A(_1031_), .Y(_740_) );
INVX2 INVX1_159_s_s_s ( .A(_879_), .Y(_754_) );
INVX2 INVX1_160_s_s_s ( .A(_1013_), .Y(_773_) );
INVX2 INVX1_161_s_s_s ( .A(_775_), .Y(_778_) );
INVX2 INVX1_162_s_s_s ( .A(_1028_), .Y(_785_) );
BUFX4 BUFX2_17_s ( .A(_1439__0_), .Y(AB[0]) );
BUFX4 BUFX2_18_s ( .A(_1439__1_), .Y(AB[1]) );
BUFX4 BUFX2_19_s ( .A(_1439__2_), .Y(AB[2]) );
BUFX4 BUFX2_20_s ( .A(_1439__3_), .Y(AB[3]) );
BUFX4 BUFX2_21_s ( .A(_1439__4_), .Y(AB[4]) );
BUFX4 BUFX2_22_s ( .A(_1439__5_), .Y(AB[5]) );
BUFX4 BUFX2_23_s ( .A(_1439__6_), .Y(AB[6]) );
BUFX4 BUFX2_24_s ( .A(_1439__7_), .Y(AB[7]) );
BUFX4 BUFX2_25_s ( .A(_1439__8_), .Y(AB[8]) );
BUFX4 BUFX2_26_s ( .A(_1439__9_), .Y(AB[9]) );
BUFX4 BUFX2_27_s ( .A(_1439__10_), .Y(AB[10]) );
BUFX4 BUFX2_28_s ( .A(_1439__11_), .Y(AB[11]) );
BUFX4 BUFX2_29_s ( .A(_1439__12_), .Y(AB[12]) );
BUFX4 BUFX2_30_s ( .A(_1439__13_), .Y(AB[13]) );
BUFX4 BUFX2_31_s ( .A(_1439__14_), .Y(AB[14]) );
BUFX4 BUFX2_32_s ( .A(_1439__15_), .Y(AB[15]) );
BUFX4 BUFX2_33_s ( .A(_1440__0_), .Y(DO[0]) );
BUFX4 BUFX2_34_s ( .A(_1440__1_), .Y(DO[1]) );
BUFX4 BUFX2_35_s ( .A(_1440__2_), .Y(DO[2]) );
BUFX4 BUFX2_36_s ( .A(_1440__3_), .Y(DO[3]) );
BUFX4 BUFX2_37_s ( .A(_1440__4_), .Y(DO[4]) );
BUFX4 BUFX2_38_s ( .A(_1440__5_), .Y(DO[5]) );
BUFX4 BUFX2_39_s ( .A(_1440__6_), .Y(DO[6]) );
BUFX4 BUFX2_40_s ( .A(_1440__7_), .Y(DO[7]) );
BUFX4 BUFX2_41_s ( .A(_1441_), .Y(WE) );
INVX4 INVX2_45_s_s_s ( .A(alu_op_3_), .Y(_1633_) );
INVX2 INVX1_163_s_s_s ( .A(alu_op_0_), .Y(_1635_) );
INVX2 INVX1_164_s_s_s ( .A(BI_5_), .Y(_1637_) );
INVX4 INVX4_8_s_s ( .A(alu_op_1_), .Y(_1639_) );
INVX2 INVX1_165_s_s_s ( .A(AI_5_), .Y(_1640_) );
INVX2 INVX1_166_s_s_s ( .A(_1638_), .Y(_1643_) );
INVX2 INVX1_167_s_s_s ( .A(_1645_), .Y(_1646_) );
INVX2 INVX1_168_s_s_s ( .A(alu_op_2_), .Y(_1647_) );
INVX2 INVX1_169_s_s_s ( .A(_1650_), .Y(_1651_) );
INVX2 INVX1_170_s_s_s ( .A(_1652_), .Y(_1653_) );
INVX4 INVX2_46_s_s_s ( .A(alu_shift_right), .Y(_1654_) );
INVX2 INVX1_171_s_s_s ( .A(_1662_), .Y(_1663_) );
INVX2 INVX1_172_s_s_s ( .A(AI_3_), .Y(_1665_) );
INVX2 INVX1_173_s_s_s ( .A(BI_2_), .Y(_1666_) );
INVX2 INVX1_174_s_s_s ( .A(AI_2_), .Y(_1668_) );
INVX1 INVX1_175_s_s ( .A(AI_1_), .Y(_1459_) );
INVX2 INVX1_176_s_s_s ( .A(BI_1_), .Y(_1460_) );
INVX2 INVX1_177_s_s_s ( .A(_1465_), .Y(_1466_) );
INVX2 INVX1_178_s_s_s ( .A(AI_0_), .Y(_1472_) );
INVX2 INVX1_179_s_s_s ( .A(BI_0_), .Y(_1473_) );
INVX2 INVX1_180_s_s_s ( .A(BI_3_), .Y(_1494_) );
INVX2 INVX1_181_s_s_s ( .A(ALU_BCD), .Y(_1506_) );
INVX2 INVX1_182_s_s_s ( .A(_1478_), .Y(_1507_) );
INVX2 INVX1_183_s_s_s ( .A(_1481_), .Y(_1509_) );
INVX2 INVX1_184_s_s_s ( .A(_1455_), .Y(_1519_) );
INVX2 INVX1_185_s_s_s ( .A(_1529_), .Y(_1530_) );
INVX2 INVX1_186_s_s_s ( .A(BI_7_), .Y(_1532_) );
INVX2 INVX1_187_s_s_s ( .A(AI_7_), .Y(_1534_) );
INVX2 INVX1_188_s_s_s ( .A(_1533_), .Y(_1537_) );
INVX2 INVX1_189_s_s_s ( .A(_1539_), .Y(_1540_) );
INVX2 INVX1_190_s_s_s ( .A(_1542_), .Y(_1543_) );
INVX2 INVX1_191_s_s_s ( .A(_1544_), .Y(_1545_) );
INVX2 INVX1_192_s_s_s ( .A(BI_6_), .Y(_1546_) );
INVX2 INVX1_193_s_s_s ( .A(AI_6_), .Y(_1548_) );
INVX2 INVX1_194_s_s_s ( .A(_1547_), .Y(_1551_) );
INVX2 INVX1_195_s_s_s ( .A(_1553_), .Y(_1554_) );
INVX2 INVX1_196_s_s_s ( .A(_1556_), .Y(_1557_) );
INVX2 INVX1_197_s_s_s ( .A(_1558_), .Y(_1559_) );
INVX2 INVX1_198_s_s_s ( .A(_1560_), .Y(_1561_) );
INVX2 INVX1_199_s_s_s ( .A(_1563_), .Y(_1564_) );
INVX2 INVX1_200_s_s_s ( .A(_1664_), .Y(_1571_) );
INVX2 INVX1_201_s_s_s ( .A(_1525_), .Y(_1573_) );
INVX2 INVX1_202_s_s_s ( .A(_1660_), .Y(_1574_) );
INVX2 INVX1_203_s_s_s ( .A(new_wire_79), .Y(_1575_) );
INVX2 INVX1_204_s_s_s ( .A(_1527_), .Y(_1593_) );
INVX2 INVX1_205_s_s_s ( .A(_1598_), .Y(_1605_) );
INVX4 INVX4_1_clone_[46]_s_s ( .A(_847_), .Y(new_wire_46) );
INVX4 INVX4_3_clone_[55]_s_s ( .A(_1099_), .Y(new_wire_55) );
INVX4 INVX4_5_clone_[62]_s_s ( .A(new_wire_63), .Y(new_wire_62) );
endmodule
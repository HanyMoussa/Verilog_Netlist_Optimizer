module testcase1 (in, out1, out2, out3, out4, out5, out6, out7, out8, out9, out10, out11, out12 , out13, out14, out15, out16, out17, out18, out19, out20);
input in;
output out1;
output out2;
output out3;
output out4;
output out5;
output out6;
output out7;
output out8;
output out9;
output out10;
output out11;
output out12;
output out13;
output out14;
output out15;
output out16;
output out17;
output out18;
output out19;
output out20;
wire vdd = 1'b1;
wire gnd = 1'b0;
INVX1 INVX1_0 ( .A(in), .Y(w1) );
INVX1 INVX1_1 ( .A(new_wire_1), .Y(out1) );
INVX1 INVX1_2 ( .A(new_wire_1), .Y(out2) );
INVX1 INVX1_3 ( .A(new_wire_2), .Y(out3) );
INVX1 INVX1_4 ( .A(new_wire_2), .Y(out4) );
INVX1 INVX1_5 ( .A(new_wire_3), .Y(out5) );
INVX1 INVX1_6 ( .A(new_wire_3), .Y(out6) );
INVX1 INVX1_7 ( .A(new_wire_4), .Y(out7) );
INVX1 INVX1_8 ( .A(new_wire_4), .Y(out8) );
INVX1 INVX1_9 ( .A(new_wire_5), .Y(out9) );
INVX1 INVX1_10 ( .A(new_wire_5), .Y(out10) );
INVX1 INVX1_11 ( .A(new_wire_6), .Y(out11) );
INVX1 INVX1_12 ( .A(new_wire_6), .Y(out12) );
INVX1 INVX1_13 ( .A(new_wire_7), .Y(out13) );
INVX1 INVX1_14 ( .A(new_wire_7), .Y(out14) );
INVX1 INVX1_15 ( .A(new_wire_8), .Y(out15) );
INVX1 INVX1_16 ( .A(new_wire_8), .Y(out16) );
INVX1 INVX1_17 ( .A(new_wire_9), .Y(out17) );
INVX1 INVX1_18 ( .A(new_wire_9), .Y(out18) );
INVX1 INVX1_19 ( .A(new_wire_10), .Y(out19) );
INVX1 INVX1_20 ( .A(new_wire_10), .Y(out20) );
BUFX2 new_buffer_1 ( .A(new_wire_11), .Y(new_wire_1) );
BUFX2 new_buffer_2 ( .A(new_wire_11), .Y(new_wire_2) );
BUFX2 new_buffer_3 ( .A(new_wire_12), .Y(new_wire_3) );
BUFX2 new_buffer_4 ( .A(new_wire_12), .Y(new_wire_4) );
BUFX2 new_buffer_5 ( .A(new_wire_13), .Y(new_wire_5) );
BUFX2 new_buffer_6 ( .A(new_wire_13), .Y(new_wire_6) );
BUFX2 new_buffer_7 ( .A(new_wire_14), .Y(new_wire_7) );
BUFX2 new_buffer_8 ( .A(new_wire_14), .Y(new_wire_8) );
BUFX2 new_buffer_9 ( .A(new_wire_15), .Y(new_wire_9) );
BUFX2 new_buffer_10 ( .A(new_wire_15), .Y(new_wire_10) );
BUFX2 new_buffer_11 ( .A(new_wire_16), .Y(new_wire_11) );
BUFX2 new_buffer_12 ( .A(new_wire_16), .Y(new_wire_12) );
BUFX2 new_buffer_13 ( .A(new_wire_17), .Y(new_wire_13) );
BUFX2 new_buffer_14 ( .A(new_wire_17), .Y(new_wire_14) );
BUFX2 new_buffer_15 ( .A(new_wire_18), .Y(new_wire_15) );
BUFX2 new_buffer_16 ( .A(new_wire_19), .Y(new_wire_16) );
BUFX2 new_buffer_17 ( .A(new_wire_19), .Y(new_wire_17) );
BUFX2 new_buffer_18 ( .A(new_wire_20), .Y(new_wire_18) );
BUFX2 new_buffer_19 ( .A(w1), .Y(new_wire_19) );
BUFX2 new_buffer_20 ( .A(w1), .Y(new_wire_20) );
endmodule
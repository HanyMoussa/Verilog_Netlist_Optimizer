module rca4 (a, b, ci, s, co);
input ci;
output co;
input [3:0] a;
input [3:0] b;
output [3:0] s;
wire vdd = 1'b1;
wire gnd = 1'b0;
OR2X2 OR2X2_1 ( .A(ci), .B(a[0]), .Y(_5_) );
NAND2X1 NAND2X1_1 ( .A(ci), .B(a[0]), .Y(_6_) );
NAND3X1 NAND3X1_1 ( .A(_4_), .B(_6_), .C(_5_), .Y(_7_) );
NOR2X1 NOR2X1_1 ( .A(ci), .B(a[0]), .Y(_1_) );
AND2X2 AND2X2_1 ( .A(ci), .B(a[0]), .Y(_2_) );
OAI21X1 OAI21X1_1 ( .A(_1_), .B(_2_), .C(b[0]), .Y(_3_) );
NAND2X1 NAND2X1_2 ( .A(_3_), .B(_7_), .Y(fa0_s) );
OAI21X1 OAI21X1_2 ( .A(_4_), .B(_1_), .C(_6_), .Y(c1) );
OR2X2 OR2X2_2 ( .A(c1), .B(a[1]), .Y(_12_) );
NAND2X1 NAND2X1_3 ( .A(c1), .B(a[1]), .Y(_13_) );
NAND3X1 NAND3X1_2 ( .A(_11_), .B(_13_), .C(_12_), .Y(_14_) );
NOR2X1 NOR2X1_2 ( .A(new_wire_1), .B(a[1]), .Y(_8_) );
AND2X2 AND2X2_2 ( .A(new_wire_1), .B(a[1]), .Y(_9_) );
OAI21X1 OAI21X1_3 ( .A(_8_), .B(_9_), .C(b[1]), .Y(_10_) );
NAND2X1 NAND2X1_4 ( .A(_10_), .B(_14_), .Y(fa1_s) );
OAI21X1 OAI21X1_4 ( .A(_11_), .B(_8_), .C(_13_), .Y(c2) );
OR2X2 OR2X2_3 ( .A(c2), .B(a[2]), .Y(_19_) );
NAND2X1 NAND2X1_5 ( .A(c2), .B(a[2]), .Y(_20_) );
NAND3X1 NAND3X1_3 ( .A(_18_), .B(_20_), .C(_19_), .Y(_21_) );
NOR2X1 NOR2X1_3 ( .A(new_wire_2), .B(a[2]), .Y(_15_) );
AND2X2 AND2X2_3 ( .A(new_wire_2), .B(a[2]), .Y(_16_) );
OAI21X1 OAI21X1_5 ( .A(_15_), .B(_16_), .C(b[2]), .Y(_17_) );
NAND2X1 NAND2X1_6 ( .A(_17_), .B(_21_), .Y(fa2_s) );
OAI21X1 OAI21X1_6 ( .A(_18_), .B(_15_), .C(_20_), .Y(c3) );
OR2X2 OR2X2_4 ( .A(c3), .B(a[3]), .Y(_26_) );
NAND2X1 NAND2X1_7 ( .A(c3), .B(a[3]), .Y(_27_) );
NAND3X1 NAND3X1_4 ( .A(_25_), .B(_27_), .C(_26_), .Y(_28_) );
NOR2X1 NOR2X1_4 ( .A(new_wire_3), .B(a[3]), .Y(_22_) );
AND2X2 AND2X2_4 ( .A(new_wire_3), .B(a[3]), .Y(_23_) );
OAI21X1 OAI21X1_7 ( .A(_22_), .B(_23_), .C(b[3]), .Y(_24_) );
NAND2X1 NAND2X1_8 ( .A(_24_), .B(_28_), .Y(fa3_s) );
OAI21X1 OAI21X1_8 ( .A(_25_), .B(_22_), .C(_27_), .Y(_0_) );
OAI21X1 OAI21X1_2_clone_[1] ( .A(new_wire_4), .B(new_wire_6), .C(new_wire_5), .Y(new_wire_1) );
OAI21X1 OAI21X1_4_clone_[2] ( .A(new_wire_7), .B(new_wire_13), .C(new_wire_8), .Y(new_wire_2) );
OAI21X1 OAI21X1_6_clone_[3] ( .A(new_wire_14), .B(new_wire_25), .C(new_wire_15), .Y(new_wire_3) );
NAND2X1 NAND2X1_1_clone_[5] ( .A(ci), .B(a[0]), .Y(new_wire_5) );
NOR2X1 NOR2X1_1_clone_[6] ( .A(ci), .B(a[0]), .Y(new_wire_6) );
NAND2X1 NAND2X1_3_clone_[8] ( .A(new_wire_9), .B(a[1]), .Y(new_wire_8) );
OAI21X1 OAI21X1_2_clone_[9] ( .A(new_wire_10), .B(new_wire_12), .C(new_wire_11), .Y(new_wire_9) );
NAND2X1 NAND2X1_1_clone_[11] ( .A(ci), .B(a[0]), .Y(new_wire_11) );
NOR2X1 NOR2X1_1_clone_[12] ( .A(ci), .B(a[0]), .Y(new_wire_12) );
NOR2X1 NOR2X1_2_clone_[13] ( .A(new_wire_24), .B(a[1]), .Y(new_wire_13) );
NAND2X1 NAND2X1_5_clone_[15] ( .A(new_wire_16), .B(a[2]), .Y(new_wire_15) );
OAI21X1 OAI21X1_4_clone_[16] ( .A(new_wire_17), .B(new_wire_23), .C(new_wire_18), .Y(new_wire_16) );
NAND2X1 NAND2X1_3_clone_[18] ( .A(new_wire_19), .B(a[1]), .Y(new_wire_18) );
OAI21X1 OAI21X1_2_clone_[19] ( .A(new_wire_20), .B(new_wire_22), .C(new_wire_21), .Y(new_wire_19) );
NAND2X1 NAND2X1_1_clone_[21] ( .A(ci), .B(a[0]), .Y(new_wire_21) );
NOR2X1 NOR2X1_1_clone_[22] ( .A(ci), .B(a[0]), .Y(new_wire_22) );
NOR2X1 NOR2X1_2_clone_[23] ( .A(new_wire_24), .B(a[1]), .Y(new_wire_23) );
OAI21X1 OAI21X1_2_clone_[1]_clone_[24] ( .A(new_wire_4), .B(new_wire_6), .C(new_wire_5), .Y(new_wire_24) );
NOR2X1 NOR2X1_3_clone_[25] ( .A(new_wire_26), .B(a[2]), .Y(new_wire_25) );
OAI21X1 OAI21X1_4_clone_[2]_clone_[26] ( .A(new_wire_7), .B(new_wire_13), .C(new_wire_8), .Y(new_wire_26) );
BUFX4 BUFX2_1_s ( .A(fa0_s), .Y(s[0]) );
BUFX4 BUFX2_2_s ( .A(fa1_s), .Y(s[1]) );
BUFX4 BUFX2_3_s ( .A(fa2_s), .Y(s[2]) );
BUFX4 BUFX2_4_s ( .A(fa3_s), .Y(s[3]) );
BUFX4 BUFX2_5_s ( .A(_0_), .Y(co) );
INVX8 INVX1_1_s_s_s ( .A(b[0]), .Y(_4_) );
INVX8 INVX1_2_s_s_s ( .A(b[1]), .Y(_11_) );
INVX8 INVX1_3_s_s_s ( .A(b[2]), .Y(_18_) );
INVX8 INVX1_4_s_s_s ( .A(b[3]), .Y(_25_) );
INVX8 INVX1_1_clone_[4]_s_s_s ( .A(b[0]), .Y(new_wire_4) );
INVX8 INVX1_2_clone_[7]_s_s_s ( .A(b[1]), .Y(new_wire_7) );
INVX8 INVX1_1_clone_[10]_s_s_s ( .A(b[0]), .Y(new_wire_10) );
INVX8 INVX1_3_clone_[14]_s_s_s ( .A(b[2]), .Y(new_wire_14) );
INVX8 INVX1_2_clone_[17]_s_s_s ( .A(b[1]), .Y(new_wire_17) );
INVX8 INVX1_1_clone_[20]_s_s_s ( .A(b[0]), .Y(new_wire_20) );
endmodule